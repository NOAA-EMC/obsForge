netcdf tms_rad_1 {
dimensions:
	spots = 11 ;
	scans = 9 ;
	channels = 12 ;
	cal_spots = 10 ;
	sensors = 6 ;
	coord = 3 ;
	coord2 = 4 ;
variables:
	float AttitudeErrorDeg(spots, scans) ;
		AttitudeErrorDeg:_FillValue = -999.f ;
		AttitudeErrorDeg:long_name = "Estimated Attitude Error" ;
		AttitudeErrorDeg:Description = "Estimated star tracker attitude error magnitude" ;
		AttitudeErrorDeg:units = "deg" ;
		AttitudeErrorDeg:Valid\ Range = 0.f, 180.f ;
	ubyte Day(scans) ;
		Day:_FillValue = 255UB ;
		Day:long_name = "UTC day" ;
		Day:Description = "UTC day of month for the nadir ADC spot." ;
		Day:units = "days" ;
		Day:Valid\ Range = 1UB, 31UB ;
	ubyte Hour(scans) ;
		Hour:_FillValue = 255UB ;
		Hour:long_name = "UTC hour" ;
		Hour:Description = "UTC hour of day for the nadir ADC spot." ;
		Hour:units = "months" ;
		Hour:Valid\ Range = 0UB, 23UB ;
	ushort Millisecond(scans) ;
		Millisecond:_FillValue = 65535US ;
		Millisecond:long_name = "UTC millisecond" ;
		Millisecond:Description = "UTC millisecond of second for the nadir ADC spot." ;
		Millisecond:units = "milliseconds" ;
		Millisecond:Valid\ Range = 0US, 999US ;
	ubyte Minute(scans) ;
		Minute:_FillValue = 255UB ;
		Minute:long_name = "UTC minute" ;
		Minute:Description = "UTC minute of our for the nadir spot." ;
		Minute:units = "minutes" ;
		Minute:Valid\ Range = 0UB, 59UB ;
	ubyte Month(scans) ;
		Month:_FillValue = 255UB ;
		Month:long_name = "UTC month" ;
		Month:Description = "UTC month of year for the nadir ADC spot." ;
		Month:units = "months" ;
		Month:Valid\ Range = 1UB, 12UB ;
	float NEDT_DS(scans, channels) ;
		NEDT_DS:_FillValue = -999.f ;
		NEDT_DS:long_name = "NEDT of cold cal. measurement" ;
		NEDT_DS:units = "K" ;
		NEDT_DS:Valid\ Range = 0.f, 100.f ;
		NEDT_DS:Description = "Estimated  NEDT  using ten samples of deep space.  Used the product of gain  (K/DN),  sample standard deviation  (DN), and normal distribution bias correction (N=10)" ;
	float NEDT_ICT(scans, channels) ;
		NEDT_ICT:_FillValue = -999.f ;
		NEDT_ICT:long_name = "NEDT of internal cal target measurement" ;
		NEDT_ICT:Description = "Estimated NEDT using ten samples viewing the internal calibration target. Used the product of gain (K/DN), sample standard deviation (DN), and normal distribution bias correction (N=10)" ;
		NEDT_ICT:units = "K" ;
		NEDT_ICT:Valid\ Range = 0.f, 100.f ;
	float NEDT_ND(scans, channels) ;
		NEDT_ND:_FillValue = -999.f ;
		NEDT_ND:long_name = "NEDT of hot cal. measurement" ;
		NEDT_ND:Description = "Estimated NEDT using ten samples with noise diode turned on viewing deep space. Used the product of gain (K/DN), sample standard deviation (DN), and normal distribution bias correction (N=10)" ;
		NEDT_ND:units = "K" ;
		NEDT_ND:Valid\ Range = 0.f, 100.f ;
	ubyte NumGPSSats(spots, scans) ;
		NumGPSSats:_FillValue = 255UB ;
		NumGPSSats:long_name = "Number of GPS satellites" ;
		NumGPSSats:Description = "Number of GPS satellites utilized for position calculation." ;
		NumGPSSats:units = "unitless" ;
		NumGPSSats:Valid\ Range = 0UB, 99UB ;
	ubyte Second(scans) ;
		Second:_FillValue = 255UB ;
		Second:long_name = "UTC second" ;
		Second:Description = "UTC second of minute for the nadir ADC spot." ;
		Second:units = "seconds" ;
		Second:Valid\ Range = 0UB, 60UB ;
	ubyte StarTrackerStatus(spots, scans) ;
		StarTrackerStatus:_FillValue = 255UB ;
		StarTrackerStatus:long_name = "Star Tracker Attitude Status Flag" ;
		StarTrackerStatus:Description = "Star Tracker Attitude Status (0=OK,1=Pending,2=Bad,3=Too_Few_Stars)" ;
		StarTrackerStatus:units = "unitless" ;
		StarTrackerStatus:Valid\ Range = 0UB, 25UB ;
	float Ta_ICT(scans, channels) ;
		Ta_ICT:_FillValue = -999.f ;
		Ta_ICT:long_name = "antenna temperature of internal cal target" ;
		Ta_ICT:units = "K" ;
		Ta_ICT:Valid\ Range = 0.f, 400.f ;
		Ta_ICT:Description = "Measured antenna temperature of the internal  calibration target, using the  noise diode as warm  cal source." ;
	ushort Year(scans) ;
		Year:_FillValue = 65535US ;
		Year:long_name = "UTC year" ;
		Year:Description = "UTC year of the nadir ADC spot." ;
		Year:units = "years" ;
		Year:Valid\ Range = 2020US, 2035US ;
	float brightness_temperature(spots, scans, channels) ;
		brightness_temperature:_FillValue = -999.f ;
		brightness_temperature:least_significant_digit = 2LL ;
		brightness_temperature:long_name = "Earth radiometric brightness temperature" ;
		brightness_temperature:units = "K" ;
		brightness_temperature:Valid\ Range = 0.f, 350.f ;
		brightness_temperature:Description = "Planck blackbody equivalent brightness temperatures  resampled to the channel 10  (G3)  boresight-Earth ellipsoid intersection." ;
	float clear_fraction(spots, scans, channels) ;
		clear_fraction:_FillValue = -999.f ;
		clear_fraction:least_significant_digit = 3LL ;
		clear_fraction:long_name = "Clear Fraction" ;
		clear_fraction:units = "Unitless" ;
		clear_fraction:Valid\ Range = 0.f, 1.f ;
		clear_fraction:Description = "Cloud-clear  fraction of each spot from time-matched geostationary satellite cloud mask, weighted by each channel\'s  antenna pattern and resampled to the channel 10  (G3) boresight-Earth ellipsoid intersection." ;
	float cold_target_counts(scans, channels) ;
		cold_target_counts:_FillValue = 0.f ;
		cold_target_counts:long_name = "Cold target counts" ;
		cold_target_counts:Description = "Mean counts (digital number) of the cold (deep space) calibration sector" ;
	ushort combinedQualityFlag(spots, scans, channels) ;
		combinedQualityFlag:_FillValue = 65535US ;
		combinedQualityFlag:long_name = "Combined Quality Flag" ;
		combinedQualityFlag:Description = "Bit 1: reserved, Bit2: non-ocean, Bit 3: Outlier timestamp, Bit 4: RFI, Bit 5: ICT-ND consistency, Bit 6: Attitude Quality, Bit 7: flagICTCal, Bit 8: flagNDCal, Bit 9: flagColdCal, Bit 10: flagPLOrientation, Bit 11: flagDayNight, Bit 12: flagAscDesc, Bit 13: flagManeuver, Bit 14: flagSolarIntrusion, Bit 15: flagLunarIntrusion" ;
		combinedQualityFlag:units = "unitless" ;
		combinedQualityFlag:Valid\ Range = 0US, 65534US ;
	float elevation(spots, scans, channels) ;
		elevation:_FillValue = -9999.f ;
		elevation:least_significant_digit = 1LL ;
		elevation:long_name = "Surface elevation" ;
		elevation:Description = "Surface elevation weighted by each channel\'s antenna pattern" ;
		elevation:units = "m" ;
		elevation:Valid\ Range = -1000.f, 10000.f ;
	ubyte flagAscDesc(spots, scans, channels) ;
		flagAscDesc:_FillValue = 255UB ;
		flagAscDesc:long_name = "Ascending/Descending flag" ;
		flagAscDesc:Description = "1 if in descending portion of orbit, 0 if in ascending portion of orbit." ;
		flagAscDesc:units = "unitless" ;
		flagAscDesc:Valid\ Range = 0UB, 1UB ;
	ubyte flagColdCal(cal_spots, scans, channels) ;
		flagColdCal:_FillValue = 255UB ;
		flagColdCal:long_name = "Cold Calibration Spot Flag" ;
		flagColdCal:Description = "Outlier detection flag for deep space calibration spots." ;
		flagColdCal:units = "unitless" ;
		flagColdCal:Valid\ Range = 0UB, 1UB ;
	ubyte flagDayNight(spots, scans, channels) ;
		flagDayNight:_FillValue = 255UB ;
		flagDayNight:long_name = "Day/Night flag" ;
		flagDayNight:Description = "1 if earth is between the sun and spacecraft, 0 if spacecraft is illuminated by sun." ;
		flagDayNight:units = "unitless" ;
		flagDayNight:Valid\ Range = 0UB, 1UB ;
	ubyte flagICTCal(cal_spots, scans, channels) ;
		flagICTCal:_FillValue = 255UB ;
		flagICTCal:long_name = "Internal Calibration Target Spot Flag" ;
		flagICTCal:Description = "Outlier detection flag for internal calibration target spots." ;
		flagICTCal:units = "unitless" ;
		flagICTCal:Valid\ Range = 0UB, 1UB ;
	ubyte flagICT_ND_Consistency(spots, scans, channels) ;
		flagICT_ND_Consistency:_FillValue = 255UB ;
		flagICT_ND_Consistency:long_name = "Internal Cal Target - Noise Diode Consistency Flag" ;
		flagICT_ND_Consistency:Description = "0 = ICT and ND are consistent, 1 = ND inconsistent with ICT thermistor, 2 = antenna_temperature_ND inconsistent with antenna_temperature_ICT, 3=Both conditions true" ;
		flagICT_ND_Consistency:units = "unitless" ;
		flagICT_ND_Consistency:Valid\ Range = 0UB, 3UB ;
	ubyte flagLunarIntrusion(spots, scans, channels) ;
		flagLunarIntrusion:_FillValue = 255UB ;
		flagLunarIntrusion:long_name = "Lunar intrusion flag" ;
		flagLunarIntrusion:Description = "1 if there is a lunar intrusion into the cold space or noise diode calibration sectors, 0 indicates no intrusion." ;
		flagLunarIntrusion:units = "unitless" ;
		flagLunarIntrusion:Valid\ Range = 0UB, 1UB ;
	ubyte flagManeuver(spots, scans, channels) ;
		flagManeuver:_FillValue = 255UB ;
		flagManeuver:long_name = "Spacecraft maneuver flag" ;
		flagManeuver:units = "unitless" ;
		flagManeuver:Valid\ Range = 0UB, 1UB ;
		flagManeuver:Description = "True if the spacecraft is in an  active  maneuver." ;
	ubyte flagNDCal(cal_spots, scans, channels) ;
		flagNDCal:_FillValue = 255UB ;
		flagNDCal:long_name = "Noise Diode Calibration Spot Flag" ;
		flagNDCal:Description = "Outlier detection flag for noise diode calibration spots." ;
		flagNDCal:units = "unitless" ;
		flagNDCal:Valid\ Range = 0UB, 1UB ;
	ubyte flagNonOcean(spots, scans, channels) ;
		flagNonOcean:_FillValue = 255UB ;
		flagNonOcean:long_name = "Non-ocean Flag" ;
		flagNonOcean:Description = "0 is ocean, 1 is land, coastline, or undefined" ;
		flagNonOcean:units = "unitless" ;
		flagNonOcean:Valid\ Range = 0UB, 1UB ;
	ubyte flagOutlierTimestamp(spots, scans) ;
		flagOutlierTimestamp:_FillValue = 255UB ;
		flagOutlierTimestamp:long_name = "Outlier Timestamp flag" ;
		flagOutlierTimestamp:Description = "1 if original spot time stamp was NaN or deviates more than 10% from expected value. These timestamps are replaced with interpolated values." ;
		flagOutlierTimestamp:units = "unitless" ;
		flagOutlierTimestamp:Valid\ Range = 0UB, 1UB ;
	ubyte flagPLOrientation(spots, scans, channels) ;
		flagPLOrientation:_FillValue = 255UB ;
		flagPLOrientation:long_name = "Payload Orientation flag" ;
		flagPLOrientation:Description = "0 if spacecraft is flying payload-first, 1 if spacecraft flying payload-aft." ;
		flagPLOrientation:units = "unitless" ;
		flagPLOrientation:Valid\ Range = 0UB, 1UB ;
	ubyte flagRFI(spots, scans, channels) ;
		flagRFI:_FillValue = 255UB ;
		flagRFI:long_name = "Radio Frequency Interference Flag" ;
		flagRFI:Description = "1 when either spacecraft or ground-source RFI is detected." ;
		flagRFI:units = "unitless" ;
		flagRFI:Valid\ Range = 0UB, 1UB ;
	ubyte flagSDRTX(spots, scans) ;
		flagSDRTX:_FillValue = 255UB ;
		flagSDRTX:long_name = "Software-defined Radio Transmit Flag" ;
		flagSDRTX:Description = "1 when the software-defined radio on the TMS bus is in transmit mode." ;
		flagSDRTX:units = "unitless" ;
		flagSDRTX:Valid\ Range = 0UB, 1UB ;
	ubyte flagSolarIntrusion(spots, scans, channels) ;
		flagSolarIntrusion:_FillValue = 255UB ;
		flagSolarIntrusion:long_name = "Solar intrusion flag" ;
		flagSolarIntrusion:Description = "1 if there is a solar intrusion into the cold space or noise diode calibration sectors, 0 indicates no intrusion." ;
		flagSolarIntrusion:units = "unitless" ;
		flagSolarIntrusion:Valid\ Range = 0UB, 1UB ;
	float instrTemp(sensors, scans) ;
		instrTemp:_FillValue = -999.f ;
		instrTemp:long_name = "Average instrument temperature" ;
		instrTemp:units = "degree Celsius" ;
		instrTemp:Valid\ Range = -50.f, 50.f ;
		instrTemp:Description = "1st:  The W/F RFE temperature; 2nd:  The G-band RFE temperature, 3-6:  ICT  thermistor temperatures." ;
	float internal_cal_target_counts(scans, channels) ;
		internal_cal_target_counts:_FillValue = 0.f ;
		internal_cal_target_counts:long_name = "Internal Calibration Target counts" ;
		internal_cal_target_counts:Description = "Mean counts (digital number) of the internal calibration target sector" ;
	float land_fraction(spots, scans, channels) ;
		land_fraction:_FillValue = -999.f ;
		land_fraction:least_significant_digit = 3LL ;
		land_fraction:long_name = "Land Fraction" ;
		land_fraction:units = "Unitless" ;
		land_fraction:Valid\ Range = 0.f, 1.f ;
		land_fraction:Description = "Land fraction weighted by each  channel\'s antenna pattern, resampled to the channel  10  (G3) boresight-Earth ellipsoid intersection." ;
	float latitude(spots, scans) ;
		latitude:_FillValue = -999.f ;
		latitude:least_significant_digit = 3LL ;
		latitude:long_name = "Latitude: line-of-sight to Earth intersection" ;
		latitude:Description = "Geodetic latitude of the line-of-sight intersection point with the Earth for each spot. Negative values are South. These correspond to the middle of each spots integration period. WGS84" ;
		latitude:units = "degree_north" ;
		latitude:Valid\ Range = -90.f, 90.f ;
	float longitude(spots, scans) ;
		longitude:_FillValue = -999.f ;
		longitude:least_significant_digit = 3LL ;
		longitude:long_name = "Longitude: line-of-sight to Earth intersection" ;
		longitude:Description = "Geodetic longitude of the line-of-sight intersection point with the Earth for each spot. Negative values are West. These correspond to the middle of each spots integration period. WGS84" ;
		longitude:units = "degree_east" ;
		longitude:Valid\ Range = -180.f, 180.f ;
	float lunar_azimuth_angle(spots, scans) ;
		lunar_azimuth_angle:_FillValue = -999.f ;
		lunar_azimuth_angle:long_name = "Line-of-sight lunar azimuth angle" ;
		lunar_azimuth_angle:Description = "The angle between the local north vector at the LOS\'s earth intersection point and a vector pointing at the center of the Moon." ;
		lunar_azimuth_angle:units = "degree" ;
		lunar_azimuth_angle:Valid\ Range = 0.f, 360.f ;
	float lunar_zenith_angle(spots, scans) ;
		lunar_zenith_angle:_FillValue = -999.f ;
		lunar_zenith_angle:long_name = "Line-of-sight lunar zenith angle" ;
		lunar_zenith_angle:Description = "The angle between the local zenith at the LOS\'s earth intersection point and a vector pointing at the center of the Moon." ;
		lunar_zenith_angle:units = "degree" ;
		lunar_zenith_angle:Valid\ Range = 0.f, 180.f ;
	float noise_diode_counts(scans, channels) ;
		noise_diode_counts:_FillValue = 0.f ;
		noise_diode_counts:long_name = "Noise diode counts" ;
		noise_diode_counts:Description = "Mean counts (digital number) of the noise diode calibration sector" ;
	float scAltitude(scans) ;
		scAltitude:_FillValue = -99999.f ;
		scAltitude:long_name = "Spacecraft altitude" ;
		scAltitude:units = "km" ;
		scAltitude:Valid\ Range = 0.f, 1000.f ;
		scAltitude:Description = "The altitude of the spacecraft above the   WGS84  ellipsoid." ;
	float scLatitude(scans) ;
		scLatitude:_FillValue = -999.f ;
		scLatitude:long_name = "Spacecraft latitude" ;
		scLatitude:Description = "The latitude of the spacecraft sub-satellite point. WGS84. " ;
		scLatitude:units = "degrees_north" ;
		scLatitude:Valid\ Range = -90.f, 90.f ;
	float scLongitude(scans) ;
		scLongitude:_FillValue = -999.f ;
		scLongitude:long_name = "Spacecraft longitude" ;
		scLongitude:Description = "The longitude of the spacecraft sub-satellite point. WGS84. " ;
		scLongitude:units = "degrees_east" ;
		scLongitude:Valid\ Range = -180.f, 180.f ;
	float scPosECEF(scans, coord) ;
		scPosECEF:_FillValue = -99999.f ;
		scPosECEF:long_name = "Spacecraft ECEF position" ;
		scPosECEF:Description = "The spacecraft position in ECEF coordinate system.  The first dimension is [x,y,z]. WGS84. Uses 41st ADC spot in each scan for timestamp." ;
		scPosECEF:units = "km" ;
		scPosECEF:Valid\ Range = -10000.f, 10000.f ;
	float scQuatECEF(scans, coord2) ;
		scQuatECEF:_FillValue = -999.f ;
		scQuatECEF:long_name = "Spacecraft Body-to-ECEF quaternion" ;
		scQuatECEF:Description = "The unit length quaternion that rotates from spacecraft body coordinate system to ECEF coordinate system.  The second dimension is [i,j,k,r], where r is the scalar element of the quaternion. WGS84. Uses 41st ADC spot in each scan for timestamp." ;
		scQuatECEF:units = "norm one" ;
		scQuatECEF:Valid\ Range = -1.f, 1.f ;
	float scRollAngle(scans) ;
		scRollAngle:_FillValue = -999.f ;
		scRollAngle:long_name = "Roll angle of the spacecraft" ;
		scRollAngle:Description = "Zero degrees means the spacecraft body Z-axis is aligned with nadir in the spacecraft body XY plane" ;
		scRollAngle:units = "degrees" ;
		scRollAngle:Valid\ Range = 0.f, 360.f ;
	float scVelECEF(scans, coord) ;
		scVelECEF:_FillValue = -99999.f ;
		scVelECEF:long_name = "Spacecraft ECEF velocity" ;
		scVelECEF:Description = "The spacecraft velocity in ECEF coordinate system.  The first dimension is [x,y,z]. WGS84. Uses 41st ADC spot in each scan for timestamp." ;
		scVelECEF:units = "km/s" ;
		scVelECEF:Valid\ Range = -10.f, 10.f ;
	float sensor_azimuth_angle(spots, scans) ;
		sensor_azimuth_angle:_FillValue = -999.f ;
		sensor_azimuth_angle:long_name = "Line-of-sight azimuth angle" ;
		sensor_azimuth_angle:units = "degree" ;
		sensor_azimuth_angle:Valid\ Range = 0.f, 360.f ;
		sensor_azimuth_angle:Description = "The angle between the local north vector at the  LOS earth intersection point and the inverse  LOS vector  (a vector pointing toward the satellite from earth)." ;
	float sensor_view_angle(spots, scans) ;
		sensor_view_angle:_FillValue = -999.f ;
		sensor_view_angle:long_name = "Line-of-sight scan angle" ;
		sensor_view_angle:Description = "The scan angle between the satellite local nadir and the Line-Of-Sight (LOS) vector from radiometer aperture." ;
		sensor_view_angle:units = "degree" ;
		sensor_view_angle:Valid\ Range = -180.f, 180.f ;
	float sensor_zenith_angle(spots, scans) ;
		sensor_zenith_angle:_FillValue = -999.f ;
		sensor_zenith_angle:long_name = "Line-of-sight zenith angle" ;
		sensor_zenith_angle:Description = "The angle between the local zenith at the LOS earth intersection point and the inverse LOS vector (a vector pointing toward the satellite from earth)." ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:Valid\ Range = 0.f, 90.f ;
	float solar_azimuth_angle(spots, scans) ;
		solar_azimuth_angle:_FillValue = -999.f ;
		solar_azimuth_angle:long_name = "Line-of-sight solar azimuth angle" ;
		solar_azimuth_angle:Description = "The angle between the local north vector at the LOS\'s earth intersection point and a vector pointing at the center of the Sun." ;
		solar_azimuth_angle:units = "degree" ;
		solar_azimuth_angle:Valid\ Range = 0.f, 360.f ;
	float solar_beta_angle(scans) ;
		solar_beta_angle:_FillValue = -999.f ;
		solar_beta_angle:long_name = "Solar beta angle" ;
		solar_beta_angle:units = "degree" ;
		solar_beta_angle:Valid\ Range = -90.f, 90.f ;
		solar_beta_angle:Description = "The angle the satellite-sun  vector extends out of the orbital plane. Uses  41st  ADC  spot in each scan for timestamp." ;
	float solar_zenith_angle(spots, scans) ;
		solar_zenith_angle:_FillValue = -999.f ;
		solar_zenith_angle:long_name = "Line-of-sight solar zenith angle" ;
		solar_zenith_angle:Description = "The angle between the local zenith at the LOS\'s earth intersection point and a vector pointing at the center of the Sun." ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:Valid\ Range = 0.f, 180.f ;

// global attributes:
		:processing_stream = "NRT" ;
		:SV_ID = 2LL ;
		:PL_ID = 3LL ;
		:DataSetQuality = "Validated" ;
		:satellite_sub_identifier = 102LL ;
		:L1BR_SW_Ver = "1.0" ;
		:version = "V01-00" ;
		:CloudMaskFiles = "" ;
		:Filename = "TMS02.1B-TBR.V01-00.NRT.ST20250915-000945.ET20250915-002141.CT20250915-013123.nc" ;
		:L1B_file = "TMS02.1B-TB.V01-00.NRT.ST20250915-000945.ET20250915-002141.CT20250915-013106.nc" ;
		:create_time = "2025-09-15T01:31:23" ;
		:start_time = "2025-09-15T00:09:45" ;
		:end_time = "2025-09-15T00:21:41" ;
		:platform = "Tomorrow-S02" ;
		:collection = "TS02_L1B-TBR" ;
		:history = "Wed Jan 14 20:06:38 2026: ncks -d scans,0,,40 -d spots,0,,8 /home/Yaping.Wang/scratchda/TMS/TS02_L1B-TBR/20250915/TMS02.1B-TBR.V01-00.NRT.ST20250915-000945.ET20250915-002141.CT20250915-013123.nc tms_rad_1_thin.nc" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 AttitudeErrorDeg =
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967,
  0.007228745, 0.01329875, 0.01441311, 0.02153408, 0.01067778, 0.007623691, 
    0.006260162, 0.007682705, 0.006368967 ;

 Day = 15, 15, 15, 15, 15, 15, 15, 15, 15 ;

 Hour = 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Millisecond = 545, 545, 545, 546, 546, 545, 546, 543, 543 ;

 Minute = 9, 11, 12, 13, 15, 16, 17, 19, 20 ;

 Month = 9, 9, 9, 9, 9, 9, 9, 9, 9 ;

 NEDT_DS =
  0.920992, 0.3366385, 0.4239399, 0.3049528, 0.3624047, 0.3597871, 0.4437959, 
    0.4654736, 0.3079226, 0.3491345, 0.3089211, 0.4935495,
  1.070568, 0.2664575, 0.3234643, 0.2626447, 0.2945721, 0.4381241, 0.567705, 
    0.4324982, 0.3836251, 0.4185684, 0.3123053, 0.3993458,
  1.366039, 0.2065686, 0.3064016, 0.2776357, 0.6128023, 0.2542739, 0.7062032, 
    0.2882292, 0.2920835, 0.4234335, 0.2626397, 0.6309291,
  0.8673847, 0.2589663, 0.3223662, 0.355191, 0.5885615, 0.4000776, 0.6225873, 
    0.4957414, 0.5862398, 0.5596453, 0.3480533, 0.5970294,
  0.9547588, 0.5113009, 0.6055072, 0.1679367, 0.2849399, 0.4114421, 
    0.4342614, 0.6373246, 0.3963611, 0.6923085, 0.3093502, 0.5944951,
  1.094337, 0.4916307, 0.3247037, 0.569667, 0.4634886, 0.3884947, 0.4494789, 
    0.8374496, 0.3694993, 0.2386155, 0.2071506, 0.5182737,
  0.8955611, 0.3246345, 0.3260876, 0.339247, 0.4508347, 0.4896194, 0.719232, 
    0.3800027, 0.4919948, 0.6295276, 0.2466143, 0.3727752,
  0.6106579, 0.3177808, 0.3897181, 0.1983792, 0.3714432, 0.3494187, 
    0.4367641, 0.5063167, 0.2602676, 0.3560435, 0.205082, 0.3610026,
  1.033536, 0.3666561, 0.3190419, 0.3933122, 0.3339703, 0.2423236, 0.731793, 
    0.5878572, 0.3155045, 0.1807157, 0.2285622, 0.3854546 ;

 NEDT_ICT =
  0.8723797, 0.7414859, 0.6686862, 0.5042081, 0.4311049, 0.6397498, 0.646958, 
    0.9128218, 0.5005927, 0.4758663, 0.680209, 0.851589,
  0.6787623, 0.6627243, 0.6828891, 0.551872, 0.8172579, 0.6672254, 0.6693863, 
    1.179067, 0.562828, 0.382894, 0.3733109, 0.6602092,
  1.025013, 0.4924738, 0.4983369, 0.920514, 0.8202181, 0.8291722, 0.7534943, 
    0.8443422, 0.3124496, 0.4421641, 0.5970457, 0.6609866,
  1.023491, 0.834868, 0.9069224, 0.6749935, 0.5482437, 0.6033021, 1.233058, 
    0.9877062, 0.5706854, 0.565797, 0.326131, 0.5992522,
  1.128208, 0.592778, 0.8047834, 0.6072147, 0.5694818, 0.8238737, 0.8051289, 
    1.034275, 0.6207725, 0.7673435, 0.5999755, 0.5460385,
  1.132068, 0.5235986, 0.586638, 0.7069965, 0.5820031, 0.7167815, 1.39631, 
    1.070724, 0.6828517, 0.2590018, 0.421341, 0.7251536,
  1.258792, 0.4786821, 0.8553205, 0.6094706, 0.3439318, 0.6878296, 0.8905503, 
    1.019783, 0.4554198, 0.5247004, 0.529409, 0.6579117,
  0.8734579, 0.5926828, 0.3955326, 0.5349962, 0.6259298, 0.7492811, 
    0.7114314, 1.407042, 0.6992438, 0.3611319, 0.3664422, 0.6590631,
  1.088963, 0.566458, 0.5522524, 0.6872014, 0.3986887, 0.7977666, 0.7310394, 
    0.6142653, 0.4844615, 0.6190645, 0.3830287, 0.7498403 ;

 NEDT_ND =
  1.274279, 0.3262446, 0.6151667, 0.4220776, 0.4755389, 0.6796814, 0.7662216, 
    0.4914381, 0.3640789, 0.5875853, 0.4019339, 0.4304799,
  1.18704, 0.5548135, 0.6416985, 0.4342254, 0.6355552, 0.7470398, 0.9644621, 
    0.8363979, 0.4391606, 0.3991137, 0.4480355, 0.8432965,
  0.7487792, 0.3621649, 0.4267796, 0.5558667, 0.4592659, 0.4985804, 
    0.9434098, 0.6349277, 0.465135, 0.4524643, 0.4519516, 0.5951023,
  1.052881, 0.3948569, 0.5783638, 0.5606439, 0.6355342, 0.7775363, 1.12645, 
    0.7116619, 0.3617051, 0.4839302, 0.4588284, 0.6450961,
  0.8971979, 0.6201425, 0.9610676, 0.5818486, 0.7718626, 0.8118398, 1.11235, 
    0.681581, 0.6243675, 0.3506402, 0.3445395, 0.5730578,
  1.039635, 0.7132221, 0.4649734, 0.5066605, 0.5913637, 0.5023276, 0.7407947, 
    0.9512028, 0.3533099, 0.6227757, 0.3199242, 0.6086825,
  1.030559, 0.4953806, 0.8183406, 0.5363894, 0.6040872, 0.5631897, 0.7792304, 
    0.7743755, 0.3464062, 0.325619, 0.5138366, 0.5298568,
  1.10875, 0.3795779, 0.5402383, 0.483402, 0.4256879, 0.4055546, 0.5200642, 
    1.239793, 0.324786, 0.265442, 0.3457287, 0.433736,
  1.461972, 0.4801933, 0.3509644, 0.5228914, 0.4006461, 0.788054, 1.101619, 
    0.8735232, 0.5338752, 0.645954, 0.3555247, 0.6160949 ;

 NumGPSSats =
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Second = 46, 6, 26, 46, 6, 26, 46, 6, 26 ;

 StarTrackerStatus =
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Ta_ICT =
  285.0699, 286.5151, 287.2558, 287.0792, 287.0522, 286.4296, 286.6774, 
    286.7286, 287.6205, 284.7508, 282.1173, 272.8118,
  286.5298, 286.3683, 286.6677, 286.7669, 286.6158, 286.2121, 285.6924, 
    286.3578, 288.4482, 285.5896, 283.1844, 275.2027,
  286.2871, 286.8028, 287.5728, 287.4896, 287.3927, 287.2058, 288.0427, 
    287.1024, 288.7872, 285.1005, 283.3649, 273.4593,
  286.5164, 287.2474, 288.6579, 287.8287, 287.6819, 287.3161, 286.8885, 
    286.6382, 288.2831, 285.8139, 283.1484, 274.4328,
  286.2985, 287.4679, 288.1561, 287.5279, 287.498, 287.208, 288.1765, 
    287.6933, 289.0677, 285.8185, 283.6646, 273.5505,
  286.26, 287.7453, 288.1312, 288.1108, 287.8557, 287.9235, 288.0897, 
    287.5548, 289.1059, 285.5457, 283.5838, 274.4954,
  285.8021, 287.1526, 287.8, 287.7933, 287.7722, 287.8084, 287.382, 287.8058, 
    289.5217, 286.8224, 283.7238, 275.704,
  284.884, 286.2217, 287.2144, 286.4338, 286.2621, 286.699, 286.7715, 
    286.1382, 288.6725, 285.3107, 283.1466, 274.027,
  284.4984, 286.2777, 287.1201, 287.0144, 286.689, 287.0005, 286.7952, 
    286.7948, 286.8681, 284.8765, 282.2299, 273.0574 ;

 Year = 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025 ;

 brightness_temperature =
  197.9453, 224.7969, 222.3516, 215.6016, 207.3516, 202.7578, 204.8516, 
    223.1797, 228.4062, 236.3672, 233.2266, 221.2266,
  194.2031, 226.9375, 223.1719, 214.3359, 204.1875, 198.6172, 198.3828, 
    213.9688, 226.4688, 237.4922, 240.8828, 231.8828,
  178.6094, 211.1484, 213.4609, 210.1875, 202.5, 196.5078, 193.7891, 
    208.7188, 222.375, 222.0625, 211.8281, 205.1797,
  171.75, 213.5312, 215.7344, 212.5312, 203.2891, 196.0312, 192.1953, 
    204.5625, 228.8516, 232.0625, 218.3125, 201.9062,
  193.8125, 226.6641, 224.3516, 213.7656, 202.8672, 194.5234, 192.5938, 
    202.0156, 225.1094, 237.0391, 244.1016, 234.4062,
  226.6562, 234.2266, 226.5938, 217.0859, 204.3672, 195.2266, 189.9844, 
    202.1953, 228.0312, 239.125, 247.2188, 243.4453,
  224.3516, 236.3281, 228.2109, 217.4141, 204.9688, 196.375, 191.9922, 
    202.7578, 230.4922, 244.1172, 254.2031, 254.1562,
  241.8281, 241.5, 231.1562, 218.6328, 204.8438, 195.0625, 191.0703, 
    203.9375, 224.9297, 239.3594, 249.7344, 257.1875,
  257.3047, 248.1875, 234.9531, 221.7812, 206.9375, 196.1641, 192.6875, 
    206.3906, 241.5859, 252.4766, 264.4531, 268.9219,
  162.6406, 195.8125, 208.0938, 213.3438, 211.4609, 204.4297, 202.1953, 
    219.6953, 210.9922, 199.0234, 187.7422, 184.5625,
  157.4062, 195.6719, 207.3516, 211.2344, 207.9922, 201.8594, 196.7656, 
    211.8906, 216.375, 205.3828, 193.2578, 186.1797,
  169.2422, 194.5781, 203.7578, 208.1719, 205.3203, 199.4766, 194.1875, 
    205.7266, 213.0625, 203.3594, 193.1172, 189.4844,
  168.2109, 198.9297, 208.7188, 211.3047, 207.0781, 199.7266, 193.7109, 
    202.5156, 219.625, 210.8594, 194.9531, 186.5781,
  165.9609, 204.2734, 213.7734, 214.6328, 208.4766, 197.1094, 192.0703, 
    200.0547, 226.6406, 223.0625, 208.6562, 201.7031,
  198.2266, 220.2188, 224.9453, 221.875, 210.9219, 200.3438, 190.4062, 
    199.8828, 232.3672, 239.9453, 239.9766, 229.1484,
  247.4141, 244.7812, 238.8672, 228.5781, 214.0469, 200.75, 192.1172, 
    198.9062, 231.6562, 242.5312, 252, 256.1172,
  240.2812, 246.1562, 242.3594, 232, 216.4062, 199.6875, 191.5078, 200.9297, 
    231.3359, 247.1172, 260.8594, 262.8125,
  255, 253.2422, 247.7891, 235.1641, 218.9688, 202.2969, 195.0234, 203.8594, 
    250.3203, 261.9453, 269.0234, 272.4609,
  161.5625, 190.7734, 203.8438, 211.6953, 211.0703, 206.5156, 201.9219, 
    217.3125, 203.2422, 191.4453, 180.1719, 177.8281,
  148.8281, 185.1719, 199.7734, 208.5781, 208.9531, 203.3594, 199.1719, 
    209.2734, 208.7656, 192.2734, 175.2969, 167.75,
  172.8984, 191.8203, 200.6328, 207.0859, 206.0234, 200.6875, 196.6641, 
    204.0625, 207.6875, 197.4531, 186.7734, 183.5859,
  171.4531, 193.2734, 202.9766, 209.3828, 207.625, 201.5156, 194.7891, 
    200.375, 206.25, 193.6641, 181.7812, 176.6484,
  166.1094, 196.5625, 208.6797, 214.6016, 211.5938, 200.7734, 192.7734, 
    199.125, 216.1641, 203.3203, 188.0234, 181.8672,
  172.9688, 201.1875, 213.0859, 216.9609, 211.7109, 200.6328, 191.5469, 
    199.6641, 229.9453, 227.8672, 214.7031, 202.7422,
  240.1562, 243.6484, 239.5938, 232.8516, 219.1016, 205.1562, 191.5781, 
    197.2891, 241.5078, 250.4531, 255.9453, 256.9219,
  248.6875, 250.6562, 246.4297, 238.1953, 223.3203, 205.125, 192.2266, 
    199.9766, 235.0469, 251.3281, 263.0391, 263.4922,
  254.7656, 255.1172, 250.2344, 240.9453, 224.0703, 207.3906, 194.5859, 
    203.2578, 257.9609, 266.5, 270.4766, 271.2188,
  161.8203, 189.1953, 201.6172, 209.9297, 211.5234, 206.8125, 204.6094, 
    216.1328, 197.6797, 186.7422, 177.875, 175.3281,
  159.6641, 185.9531, 200.1484, 207.3359, 209.8281, 204.2812, 199, 209.2031, 
    202.3047, 186.2344, 170.9141, 166.0156,
  172.0391, 190.4219, 199.3906, 205.7969, 206.1719, 200.8984, 196.3281, 
    204.4141, 202.7969, 191.3906, 182.875, 178.6875,
  165.2578, 185.875, 198.7188, 205.6172, 206.9141, 201.2969, 195.0156, 
    199.8828, 199.625, 183.2031, 169.7188, 164.9297,
  167.3516, 191.8828, 204.2891, 211.0312, 211.7578, 201.0781, 194.7734, 
    198.0547, 201.4766, 188.5625, 175.5938, 171.2969,
  168.5469, 194.4219, 206.5234, 212.6562, 212.2891, 201.8281, 192.8438, 
    197.3516, 218.125, 207.4375, 197.5391, 193.8672,
  220.5, 233.0703, 235.0156, 231.6172, 221.3828, 206.0234, 193.6328, 
    196.3359, 239.5781, 248.4141, 251.2031, 240.9219,
  248.3516, 250.9531, 249.2344, 241.5859, 227.3125, 207.7266, 193.9219, 
    198.5312, 236.9688, 252.2344, 261.9219, 260.7891,
  257.6797, 256.5234, 253.7344, 244.625, 229.6094, 210.9688, 197.8516, 
    201.4766, 260.0781, 267.1406, 271.9141, 271.4531,
  160.5469, 184.7812, 197.5, 206.9609, 210.7031, 207.1172, 204.5469, 
    215.4766, 191.6719, 176.0391, 165.3672, 161.2031,
  162.6719, 184.4141, 196.3438, 205.7656, 207.9844, 204.7969, 199.1875, 
    209.1562, 198.5391, 183.7344, 171.6562, 167.5625,
  169.1797, 186.8516, 196.1641, 204.2031, 205.3047, 201.0625, 195.9062, 
    202.375, 199.8281, 189.25, 180.6719, 176.2891,
  168.2891, 186.4531, 198.2266, 204.9766, 206.5625, 201.8125, 194.2344, 
    199.3438, 198.9922, 183.9688, 171.4688, 166.1484,
  172.7031, 192.2578, 203.3516, 209.2422, 210.7266, 203.7734, 194.9844, 
    197.4922, 215.2266, 201.0391, 184.6094, 175.2656,
  168.3594, 190.6562, 202.6016, 210.4609, 212.0156, 204.2344, 193.9844, 
    196.4609, 213.9844, 201.6172, 190.6016, 187.5234,
  220.4062, 229.7734, 232.6172, 231.3516, 221.9375, 207.1641, 194.3125, 
    197.7891, 236.2109, 243.5859, 241.0078, 223.7656,
  255.2812, 252.3828, 248.9297, 241.5156, 227.9531, 209.25, 193.9453, 
    198.3672, 237.4922, 249.6953, 257.9062, 259.9609,
  257.7031, 256.9844, 253.375, 244.7109, 232.8516, 212.4297, 197.6484, 
    204.4922, 260.5078, 267.5625, 272.2266, 269.6875,
  155.8281, 181.3359, 194.3906, 205.3906, 208.8906, 206.3516, 203.7734, 
    216.4297, 189.2344, 172.9062, 162.0938, 160.0234,
  163.2891, 186.7578, 197.1641, 204.625, 206.5859, 203.9922, 201.4375, 
    208.1953, 200.0391, 187.2734, 177.9688, 174.3359,
  168.5547, 186.7578, 194.7109, 203.4688, 204.5625, 201.3047, 196.4219, 
    203.4688, 196.5, 186.2031, 178.5, 175.8516,
  172.4375, 189.8594, 199.2109, 207.0859, 207.0938, 201.2344, 194.2656, 
    199.9766, 208.9609, 196.3516, 184.125, 179.3906,
  173.8438, 192.1016, 201.8594, 209.8672, 209.2422, 203.4609, 193.4844, 
    197.9219, 217.3594, 203.6172, 185.5625, 175.9688,
  170.5547, 191.0859, 201.5625, 209.2578, 211.3828, 204.3516, 194.2422, 
    198.1172, 214.6875, 203.2422, 192.6875, 188.6484,
  216.3906, 228.3516, 231.5938, 230.6875, 222, 206.5781, 193.9453, 197.6953, 
    235.7109, 243.2188, 238.9453, 221.2188,
  247.7266, 248.1797, 246.0547, 241, 228.4609, 211.0625, 195.7188, 200.3828, 
    236.0547, 247.9219, 257.2188, 254.6875,
  252.8203, 255.1641, 253.1094, 246.1641, 231.8047, 212.7578, 198.0547, 
    203.25, 260.5938, 267.0391, 270.1172, 267.5859,
  158.75, 180.8438, 193.3672, 203.9297, 208.6406, 205.8125, 204.7578, 
    216.1484, 192.8438, 177.0703, 165.9453, 163.1875,
  161.5391, 183.5938, 194.4688, 202.6016, 206.6953, 203.9609, 198.2734, 
    210.8438, 194.0391, 181.3359, 172.0469, 169.1953,
  165.1719, 180.125, 191.2344, 200.6719, 204.2734, 201.4375, 196.4219, 
    203.4688, 189.4688, 176.6562, 168.7578, 165.5391,
  169.7812, 188.4766, 198.8594, 205.8984, 206.9844, 201.25, 194.4922, 
    201.0312, 210.9609, 196.8594, 181.6953, 177.8281,
  171.5156, 190.9453, 201.0078, 208.3594, 208.3516, 202.1094, 193.3984, 
    198.9453, 214.6797, 200.8984, 187.1562, 178.375,
  173.1641, 192.7109, 202.6719, 209.5859, 210.875, 203.3516, 193.8359, 
    198.3594, 209.9922, 199.3984, 191.0391, 187.8125,
  216.5469, 228.7344, 232.3281, 230.3203, 222.0781, 206.3984, 193.2188, 
    198.3438, 239.4453, 245.9141, 236.7344, 220.1953,
  236.2891, 242.3828, 242.9062, 238.0391, 227.9062, 210.4219, 194.8906, 
    200.625, 235.9922, 246.5469, 249.9141, 241.9609,
  255.1406, 254.75, 252.4375, 245.0938, 230.9141, 213.2031, 198.9453, 
    205.1875, 260.625, 266.5859, 269.7344, 268.9375,
  156.2578, 179.9688, 195.4609, 204.9922, 208.4297, 206.5078, 202.8672, 
    218.4453, 195.9922, 180.8828, 168.8906, 166.2188,
  155.7734, 179.7656, 191.8906, 201.9688, 206.3359, 203.3281, 199.1328, 
    210.7266, 189.4453, 175.7891, 165.8594, 163.1719,
  160.5781, 178.5, 190.4141, 199.1875, 203.2656, 199.9922, 195.5703, 
    205.5391, 186.7109, 173.2266, 164.2734, 162.6719,
  162.3359, 181.5547, 193.1953, 201.9688, 204.9219, 199.75, 193.5859, 
    200.875, 206.1484, 190.0234, 173.8359, 167.3125,
  167.25, 188.4766, 198.9453, 207.1016, 206.5703, 200.2578, 193.8359, 
    197.4375, 216.7734, 203.5625, 189, 182.0312,
  179.8438, 194.9062, 204.5156, 210.9766, 209.7891, 202.6016, 193.6562, 
    200.6016, 214.9297, 205.2188, 198.0312, 195.8438,
  228.1406, 234.6016, 236.6875, 233.1953, 221.6328, 205.6484, 194.1484, 
    198.4609, 242.6172, 249.4688, 242.9375, 225.7188,
  236.0547, 240.25, 240.9219, 238.2578, 225.7969, 208.8281, 195.8594, 
    200.5781, 237.2812, 248.7266, 251.5, 238.1484,
  244.5625, 249.2188, 249.2266, 241.2188, 228.4375, 210.6484, 200.2578, 
    206.2656, 250.3906, 260.8203, 266.25, 264.0312,
  161.5703, 186.3594, 199.6094, 208.4062, 208.6484, 204.6562, 203.7188, 
    219.2812, 201.3047, 188.6094, 178.4844, 175.6641,
  154.9375, 180.8125, 193.625, 202.9531, 205.2578, 202.5078, 199.4062, 
    213.8281, 192.8203, 178.3359, 167.6172, 165.8281,
  168.6016, 187.4062, 198.9297, 205.8203, 206.1172, 199.1562, 195.2578, 
    207.2578, 195.0547, 183.7109, 175.1328, 172.0859,
  158.7188, 182.0703, 195.2578, 203.3359, 204.4688, 197.5156, 192.3984, 
    203.9688, 208.5781, 189.4141, 168.5781, 160.75,
  167.1797, 189.5859, 200.0625, 205.8672, 205.9453, 198.9141, 192.4766, 
    201.8047, 212.1094, 199.4844, 188.0547, 183.0547,
  191.5781, 207.5391, 212.8359, 214.7344, 209.9219, 201.4453, 192.7344, 
    197.75, 224.0078, 217.2969, 209.9688, 206.9688,
  227, 234.7266, 235.8594, 230.1484, 216.9609, 203.6094, 191.8047, 200.2266, 
    244.3984, 250.6719, 246.2812, 232.5938,
  232.7578, 239.1719, 240.0312, 234.7656, 222.9609, 206.4844, 195.0703, 
    203.0391, 236.8359, 249.6484, 249.0625, 236.0547,
  241.8984, 245.8203, 245.1719, 239.0156, 224.5859, 209.0156, 199.9531, 
    208.9766, 238.0625, 249.2188, 258.75, 259.6562,
  165.8359, 194.2031, 206.4453, 211.5, 209.7656, 204.4141, 203.7891, 
    224.6094, 205.2266, 194.3516, 186.1016, 182.6406,
  158.1484, 184.8438, 196.2734, 204.6328, 204.6016, 201.8047, 198.9609, 
    217.1016, 200.9297, 187.3125, 174.9219, 170.2188,
  168.5625, 196.0078, 205.4844, 208.8203, 204.2812, 197.1328, 193.125, 
    211.1797, 204.6953, 197.1406, 191.7969, 188.8203,
  162.5703, 191.5078, 202.6641, 207.0469, 204.1328, 196.0312, 192.2109, 
    205.875, 211.6953, 197.1016, 179.5469, 172.1797,
  180.4688, 201.4688, 209.5234, 211.0547, 205.8672, 196.8594, 192.1406, 
    205.7422, 220.5, 212.3828, 203.7344, 199.2891,
  204.4922, 222.0469, 224.3203, 219.6016, 208.0391, 198.7188, 192.0625, 
    201.7812, 237.1406, 240.9922, 233.2891, 223.1328,
  219.5703, 232.2422, 231.4297, 224.9062, 211.9062, 201.3203, 193.8438, 
    202.7109, 241.1484, 249.3594, 250.9062, 239.5625,
  228.6953, 238.6406, 237.6875, 229.0859, 217.4609, 202.375, 197.9062, 
    207.6953, 244.5312, 253.0547, 251.4844, 238.5781,
  217.9141, 236.2266, 238.7891, 232.2812, 219.6641, 206.0312, 200.0391, 
    212.0156, 238.3359, 248.7422, 251.8516, 238.8438,
  171.8984, 210.2734, 215.1641, 213.0781, 208.6172, 205.8281, 211.8047, 
    232.7109, 220.7656, 214.7266, 200.3281, 191.4297,
  174.9375, 203.3203, 209.6953, 209.8047, 204.4531, 200.9609, 202.0938, 
    225.8047, 215.5156, 206.2031, 191.6328, 184.1484,
  166.3125, 211.0234, 215.6406, 211.7422, 201.8984, 195.5234, 197, 221.1328, 
    224.4453, 216.2891, 205.7891, 196.625,
  166.875, 205.1328, 210.9062, 208.0859, 199.9297, 192.6953, 194.6406, 
    214.3672, 218.4453, 205.8203, 189.5547, 181.8438,
  190.6953, 216.7734, 218.0156, 211.5703, 201.5547, 193.2188, 194.1016, 
    211.9531, 225.2734, 226.9141, 218, 209.9375,
  227.9062, 231.4297, 223.3203, 213.1016, 202.6641, 196.7656, 193.4688, 
    210.6562, 230.6641, 240.6016, 248.0547, 241.6406,
  213.5703, 228.7734, 224.2109, 215.2109, 205.4219, 198.7188, 197.0234, 
    213.4375, 230.8203, 240.5625, 244.9922, 231.4141,
  219.0234, 232.9688, 228.6172, 219.8203, 210.7891, 202.9062, 202.4062, 
    216.3203, 239.875, 247.7188, 248.7422, 238.5469,
  216.0312, 235.7031, 231.6172, 224.1484, 214.6797, 207.7656, 208.2812, 
    220.1328, 246.6406, 251.8828, 249.8828, 236.9297 ;

 clear_fraction =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 cold_target_counts =
  -135331, 5.215981e+10, 2.747025e+10, 8.766734e+10, 6.284173e+10, 
    6.886358e+10, 1.638252e+10, 1.825988e+10, -401073, -305549.6, -248527.8, 
    -369292,
  -135447.2, 5.210318e+10, 2.748089e+10, 8.770406e+10, 6.279555e+10, 
    6.878152e+10, 1.637369e+10, 1.82421e+10, -401024.3, -306055.1, -248482, 
    -369764.8,
  -135388.2, 5.222802e+10, 2.751996e+10, 8.781498e+10, 6.295732e+10, 
    6.899217e+10, 1.641618e+10, 1.829135e+10, -401167.5, -305505, -248567.4, 
    -369701.4,
  -135227, 5.226679e+10, 2.753038e+10, 8.784935e+10, 6.293148e+10, 
    6.897811e+10, 1.641695e+10, 1.830196e+10, -401277.7, -305750.7, 
    -247987.1, -369341.3,
  -135267.5, 5.23825e+10, 2.759822e+10, 8.808477e+10, 6.315346e+10, 
    6.916601e+10, 1.644827e+10, 1.834374e+10, -400146.2, -305171.2, 
    -247617.1, -368432.9,
  -135177.5, 5.241857e+10, 2.759802e+10, 8.807775e+10, 6.311945e+10, 
    6.914515e+10, 1.645951e+10, 1.833085e+10, -400248.8, -305150.4, 
    -247751.5, -368547.3,
  -135432.9, 5.240149e+10, 2.760304e+10, 8.806408e+10, 6.309915e+10, 
    6.914725e+10, 1.645113e+10, 1.835318e+10, -400292.1, -305282.1, 
    -247842.5, -368195.4,
  -135069.6, 5.24199e+10, 2.758828e+10, 8.804146e+10, 6.309356e+10, 
    6.916003e+10, 1.645017e+10, 1.831321e+10, -399356.1, -304548.7, 
    -247282.3, -367910.6,
  -134302.8, 5.257093e+10, 2.765796e+10, 8.828454e+10, 6.318433e+10, 
    6.921183e+10, 1.647122e+10, 1.834723e+10, -398754.3, -304431.3, -247111, 
    -366712.5 ;

 combinedQualityFlag =
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2306,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2306,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2306,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2322,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2322,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2322,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2322,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026, 1026,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2322,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2322,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2306,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2066,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 18,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2306,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050, 2050,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 258, 2,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024,
  1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024, 1024 ;

 elevation =
  119.25, 111.8125, 117.6875, 113.3125, 115, 115.875, 115, 114.625, 55.9375, 
    54.8125, 56.5, 54.75,
  85.75, 89.0625, 82.25, 87.6875, 89.125, 89.25, 89, 88.875, 63, 63, 63, 
    61.875,
  2417.438, 2497.5, 2481.25, 2493.625, 2493.188, 2493.438, 2493.438, 
    2492.688, 2416.875, 2414.625, 2416.5, 2415.875,
  1914.25, 1958.25, 1944.812, 1954.5, 1955.312, 1956.062, 1954.938, 1954.438, 
    1959.062, 1961.812, 1958.812, 1959.688,
  666.0625, 706.75, 689.625, 701.9375, 703.9375, 705.3125, 702.625, 701.5625, 
    687.9375, 680.375, 690.6875, 689.75,
  155.8125, 143.125, 140.8125, 144.25, 146.3125, 147.125, 145.1875, 144.25, 
    50.5, 46.125, 46.4375, 44.6875,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2414.5, 2418.938, 2417.188, 2418.375, 2418.75, 2418.875, 2418.5, 2418.375, 
    2420.188, 2420.375, 2420.688, 2420.562,
  2390.812, 2392.375, 2391.75, 2392.125, 2392, 2391.875, 2392.188, 2392.25, 
    2387.812, 2387.875, 2388.125, 2387.75,
  3124.75, 3127.312, 3126.625, 3127.062, 3127, 3127, 3127.062, 3127.062, 
    3127.125, 3127, 3127.375, 3127.375,
  2710.812, 2714.062, 2713, 2713.812, 2713.875, 2714, 2713.812, 2713.75, 
    2713.5, 2713.125, 2713.625, 2713.688,
  1945.062, 1943.562, 1943.062, 1943.375, 1943.938, 1944.125, 1943.5, 
    1943.375, 1945.188, 1945, 1944.938, 1945.062,
  1839.375, 1858.375, 1850.5, 1855.625, 1856.625, 1857.5, 1856, 1855.562, 
    1868.125, 1866.688, 1870, 1870.125,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2593.938, 2596.875, 2595.875, 2596.562, 2596.625, 2596.688, 2596.625, 
    2596.562, 2595.75, 2595.875, 2595.938, 2595.875,
  2766.188, 2769.75, 2768.75, 2769.438, 2769.312, 2769.25, 2769.375, 
    2769.375, 2766.688, 2766.562, 2766.938, 2766.812,
  3250.688, 3254.875, 3253.812, 3254.562, 3254.562, 3254.562, 3254.625, 
    3254.562, 3250.312, 3250.062, 3250.312, 3250.188,
  2907, 2908.75, 2907.438, 2908.312, 2908.75, 2909, 2908.438, 2908.25, 
    2908.562, 2908.062, 2908.438, 2908.562,
  2419.688, 2427.375, 2424.688, 2426.5, 2426.688, 2426.75, 2426.562, 2426.5, 
    2424.688, 2424.062, 2425.125, 2425.062,
  2416.562, 2420.688, 2418.938, 2420.125, 2420.125, 2420.125, 2420.188, 
    2420.125, 2418.875, 2418.438, 2419.25, 2419.062,
  172.125, 204.8125, 192.9375, 200.1875, 200.375, 200.5, 199.8125, 199.8125, 
    246.5625, 245.4375, 251, 250.4375,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2784.375, 2786.125, 2785.375, 2785.875, 2786.062, 2786.188, 2786, 2785.938, 
    2785.5, 2785.562, 2785.625, 2785.5,
  3007.688, 3011.312, 3010.25, 3010.938, 3010.875, 3010.875, 3011, 3010.938, 
    3008.562, 3008.312, 3008.75, 3008.625,
  3450.188, 3453.25, 3452.375, 3452.938, 3452.938, 3452.875, 3453, 3452.938, 
    3450.812, 3450.688, 3450.938, 3450.875,
  3213.062, 3214.562, 3213.625, 3214.312, 3214.75, 3215, 3214.5, 3214.375, 
    3214.125, 3213.688, 3214.062, 3214.312,
  2766.312, 2769.875, 2768.438, 2769.5, 2769.438, 2769.5, 2769.5, 2769.438, 
    2765.25, 2764.875, 2765.312, 2765.25,
  2716, 2719.75, 2718.375, 2719.375, 2719.5, 2719.5, 2719.375, 2719.312, 
    2716.625, 2716.312, 2716.875, 2716.812,
  122.75, 116.5, 117.6875, 117.0625, 117.25, 117.375, 117.25, 117, 84.9375, 
    84.125, 83.125, 82.5625,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2981, 2984.062, 2982.938, 2983.688, 2983.812, 2983.812, 2983.75, 2983.688, 
    2982.625, 2982.75, 2982.375, 2982.5,
  3187.125, 3189.562, 3188.875, 3189.312, 3189.25, 3189.25, 3189.312, 
    3189.312, 3188.188, 3188.062, 3188.438, 3188.375,
  3616.375, 3619, 3618.25, 3618.812, 3618.75, 3618.75, 3618.812, 3618.812, 
    3616.25, 3616.125, 3616.562, 3616.562,
  3417.188, 3418.25, 3417.75, 3418.188, 3418.438, 3418.562, 3418.125, 
    3418.062, 3416.688, 3416.375, 3416.562, 3416.625,
  3017.062, 3019.812, 3018.938, 3019.5, 3019.625, 3019.688, 3019.562, 3019.5, 
    3017.312, 3016.938, 3017.25, 3017.25,
  2970.312, 2972.312, 2971.375, 2972.062, 2972.188, 2972.25, 2972.062, 2972, 
    2971.312, 2971, 2971.375, 2971.375,
  71.625, 71.4375, 71.3125, 71.3125, 71.4375, 71.4375, 71.3125, 71.3125, 
    72.9375, 73, 73, 72.9375,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3170.312, 3172.688, 3171.875, 3172.5, 3172.375, 3172.375, 3172.5, 3172.438, 
    3171.875, 3172, 3171.75, 3171.75,
  3306.938, 3307.75, 3307.5, 3307.688, 3307.625, 3307.625, 3307.75, 3307.75, 
    3305.5, 3305.438, 3305.5, 3305.438,
  3785.812, 3788.875, 3788, 3788.75, 3788.625, 3788.625, 3788.625, 3788.625, 
    3786.125, 3785.875, 3786.312, 3786.125,
  3563.562, 3563.875, 3563.688, 3563.938, 3564.062, 3564.125, 3563.938, 
    3563.875, 3562.562, 3562.438, 3562.438, 3562.5,
  3222.938, 3225.688, 3224.688, 3225.438, 3225.562, 3225.625, 3225.438, 
    3225.438, 3224.5, 3224.062, 3224.625, 3224.5,
  3140.875, 3142.688, 3141.812, 3142.312, 3142.5, 3142.625, 3142.375, 
    3142.312, 3143.812, 3143.625, 3144, 3144,
  53, 52.8125, 52.875, 52.875, 52.8125, 52.8125, 52.8125, 52.8125, 54.125, 
    54.1875, 54.125, 54.1875,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3264.125, 3265.312, 3264.812, 3265.125, 3265.188, 3265.188, 3265.188, 
    3265.125, 3265.188, 3265.25, 3265.25, 3265.25,
  3408.625, 3409.875, 3409.312, 3409.812, 3409.688, 3409.688, 3409.75, 
    3409.75, 3407.688, 3407.5, 3407.75, 3407.688,
  3953.938, 3955, 3954.688, 3954.938, 3954.812, 3954.812, 3954.938, 3954.938, 
    3952.438, 3952.438, 3952.438, 3952.375,
  3704.375, 3706.062, 3705.438, 3705.812, 3706, 3706.125, 3705.938, 3705.875, 
    3704.5, 3704.188, 3704.438, 3704.375,
  3375.75, 3378.375, 3377.562, 3378.188, 3378.188, 3378.25, 3378.188, 
    3378.125, 3376.125, 3375.812, 3376.125, 3376.125,
  3280.812, 3281.688, 3281.188, 3281.5, 3281.75, 3281.812, 3281.562, 3281.5, 
    3281.875, 3281.688, 3281.938, 3281.938,
  41.1875, 40.5625, 41, 40.9375, 41.125, 41.25, 40.875, 40.8125, 39.25, 
    39.1875, 38.9375, 39.0625,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3228.875, 3227.438, 3227.938, 3227.625, 3227.625, 3227.625, 3227.562, 
    3227.625, 3228.438, 3228.438, 3228.562, 3228.562,
  3530.812, 3531.125, 3531, 3531.125, 3531.125, 3531.125, 3531.188, 3531.188, 
    3529.5, 3529.438, 3529.438, 3529.438,
  4040, 4041, 4041, 4041, 4040.875, 4040.812, 4041, 4041, 4040.188, 4040.188, 
    4040.25, 4040.25,
  3751.5, 3750.75, 3751.188, 3750.938, 3750.938, 3750.875, 3750.875, 
    3750.875, 3752.125, 3752.25, 3752.125, 3752.062,
  3542.5, 3544, 3543.375, 3543.875, 3543.938, 3544, 3543.812, 3543.812, 
    3542.312, 3542.062, 3542.438, 3542.375,
  3330.375, 3329.5, 3329.562, 3329.438, 3329.75, 3329.812, 3329.5, 3329.438, 
    3331.062, 3331, 3330.812, 3331,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3139.875, 3138.438, 3138.875, 3138.562, 3138.562, 3138.5, 3138.562, 
    3138.562, 3140.25, 3140.25, 3140.375, 3140.438,
  3595.938, 3597.938, 3597.438, 3597.688, 3597.5, 3597.375, 3597.688, 
    3597.688, 3596.938, 3596.938, 3597.25, 3597.062,
  3676.438, 3664.688, 3669.375, 3666.188, 3665.875, 3665.5, 3666, 3666.25, 
    3667.125, 3668.75, 3666.5, 3666.25,
  3586.062, 3584.25, 3585.312, 3584.5, 3584.375, 3584.312, 3584.5, 3584.562, 
    3585.5, 3585.875, 3585.5, 3585.562,
  3714.062, 3714.125, 3714.312, 3714.188, 3714.25, 3714.312, 3714.062, 
    3714.062, 3717.062, 3717.125, 3717.188, 3717.312,
  3008.312, 2999.562, 3003.125, 3000.875, 3001, 3001.062, 3000.375, 3000.438, 
    3009.562, 3010.75, 3009.438, 3009.562,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2905.438, 2903.312, 2904.625, 2903.625, 2903.5, 2903.375, 2903.562, 
    2903.688, 2906.688, 2906.75, 2906.75, 2907,
  3634.5, 3635.25, 3635.438, 3635.312, 3635, 3634.875, 3635.25, 3635.312, 
    3634.875, 3635, 3635.062, 3635,
  2945.5, 2936.438, 2939.375, 2937.25, 2937.312, 2937.312, 2937.312, 
    2937.375, 2938.938, 2939.625, 2937.812, 2938.125,
  3276.25, 3273.938, 3275.562, 3274.25, 3273.812, 3273.562, 3274.188, 
    3274.375, 3277.312, 3278.062, 3277.375, 3277.375,
  3393.375, 3385.312, 3387.812, 3385.938, 3386.125, 3386.25, 3385.938, 3386, 
    3390.625, 3391.375, 3390.188, 3390.375,
  1200.188, 1171, 1179.75, 1173.125, 1173.188, 1173.375, 1173.375, 1173.688, 
    1211.25, 1214.062, 1211.062, 1212.688,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2467.062, 2464.062, 2467.688, 2465.188, 2465.062, 2464.562, 2464.438, 
    2464.75, 2480.688, 2480.562, 2480.062, 2481.438,
  3168.562, 3154.938, 3160.75, 3156.438, 3156.25, 3155.875, 3156.312, 
    3156.688, 3175.875, 3178.75, 3175.062, 3175.875,
  2031.688, 2004.812, 2011.375, 2006.562, 2009, 2009.688, 2007.562, 2007.75, 
    2059.812, 2064.688, 2057.75, 2061.188,
  2663.938, 2673.25, 2673.188, 2674, 2670.938, 2670.375, 2672, 2672.125, 
    2667.875, 2666.812, 2668.875, 2667.75,
  2284.688, 2245.188, 2257.062, 2248.312, 2248.812, 2249.062, 2248.062, 
    2248.25, 2273.875, 2277, 2271.812, 2273.188,
  0.5, 0.125, 0.1875, 0.125, 0.125, 0.125, 0.125, 0.125, 0.0625, 0.0625, 
    0.0625, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagAscDesc =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagColdCal =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagDayNight =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 flagICTCal =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagICT_ND_Consistency =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagLunarIntrusion =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagManeuver =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagNDCal =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagNonOcean =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagOutlierTimestamp =
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagPLOrientation =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagRFI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagSDRTX =
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagSolarIntrusion =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 instrTemp =
  7.157745, 7.322113, 7.232147, 7.329926, 7.239929, 7.239929, 7.239929, 
    7.149994, 6.985718,
  4.123993, 4.117188, 4.117188, 4.041748, 3.95282, 3.870667, 3.870667, 
    3.870667, 3.706299,
  14.73795, 14.93597, 15.19318, 15.29208, 15.41064, 15.52914, 15.48969, 
    15.5687, 15.17337,
  14.63879, 14.87659, 15.07452, 15.25253, 15.41064, 15.62793, 15.9043, 
    15.78589, 15.35132,
  15.03497, 15.35132, 15.54895, 15.58844, 15.82535, 15.98325, 16.02267, 
    15.9043, 15.46991,
  13.92313, 14.12231, 14.26154, 14.51981, 14.63879, 14.75775, 15.11411, 
    15.07452, 14.75775 ;

 internal_cal_target_counts =
  -195076.2, 8.491579e+10, 4.444597e+10, 1.499882e+11, 1.077749e+11, 
    1.175158e+11, 2.806778e+10, 3.114601e+10, -540468, -401457.3, -342147.2, 
    -478669.7,
  -195573.1, 8.502474e+10, 4.44778e+10, 1.500758e+11, 1.078564e+11, 
    1.17654e+11, 2.808893e+10, 3.116933e+10, -541344.8, -402522.9, -342356.2, 
    -480145.2,
  -195640.1, 8.510062e+10, 4.453539e+10, 1.502858e+11, 1.080352e+11, 
    1.17835e+11, 2.815648e+10, 3.119877e+10, -541406.5, -402212.9, -342639.6, 
    -480068.7,
  -195631.5, 8.5159e+10, 4.458624e+10, 1.504267e+11, 1.080965e+11, 
    1.179348e+11, 2.814965e+10, 3.121333e+10, -541414.3, -401958.2, -342026, 
    -479791.3,
  -195401.6, 8.541504e+10, 4.469936e+10, 1.508563e+11, 1.083788e+11, 
    1.182063e+11, 2.821678e+10, 3.1311e+10, -540577.6, -401892, -341736.6, 
    -478867.5,
  -195390.3, 8.554936e+10, 4.474583e+10, 1.510902e+11, 1.085485e+11, 
    1.183384e+11, 2.827912e+10, 3.13555e+10, -540611.7, -401747.7, -341784.6, 
    -478786.7,
  -195411.4, 8.549841e+10, 4.472888e+10, 1.509934e+11, 1.084413e+11, 
    1.183053e+11, 2.824327e+10, 3.133146e+10, -540564.8, -401874.4, 
    -341823.9, -478963.7,
  -194598.6, 8.547795e+10, 4.470493e+10, 1.507942e+11, 1.08312e+11, 
    1.182233e+11, 2.823254e+10, 3.128787e+10, -539266.2, -400824.6, 
    -341072.7, -477997.8,
  -193652.1, 8.570545e+10, 4.478925e+10, 1.511565e+11, 1.085909e+11, 
    1.184257e+11, 2.827033e+10, 3.135478e+10, -537981.7, -400853.5, 
    -340588.4, -476046.5 ;

 land_fraction =
  0.7763672, 0.8388672, 0.8173828, 0.8310547, 0.8300781, 0.8291016, 
    0.8310547, 0.8320312, 0.9453125, 0.9501953, 0.9492188, 0.953125,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.21875, 0.2050781, 0.2001953, 0.2060547, 0.2089844, 0.2099609, 0.2080078, 
    0.2070312, 0.09082031, 0.08398438, 0.08496094, 0.08496094,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.6855469, 0.7451172, 0.7197266, 0.7373047, 0.7382812, 0.7392578, 
    0.7363281, 0.7353516, 0.8125, 0.8085938, 0.8193359, 0.8212891,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9980469, 0.9980469, 0.9970703, 0.9980469, 0.9980469, 0.9980469, 
    0.9970703, 0.9970703, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8251953, 0.8310547, 0.8212891, 0.8261719, 0.8291016, 0.8310547, 
    0.8251953, 0.8251953, 0.9570312, 0.9589844, 0.9628906, 0.9609375,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.0078125, 0.001953125, 0.002929688, 0.001953125, 0.001953125, 0.001953125, 
    0.001953125, 0.001953125, 0.0009765625, 0.0009765625, 0.0009765625, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 latitude =
  -77.8252, -82.68164, -87.0791, -86.38379, -81.78613, -76.90137, -71.97168, 
    -66.99316, -62.02539,
  -77.77637, -82.68359, -87.19141, -86.47168, -81.81055, -76.89258, 
    -71.91699, -66.93555, -61.93066,
  -77.28613, -81.91016, -85.56836, -85.0752, -81.1084, -76.42969, -71.56348, 
    -66.64355, -61.67285,
  -76.79199, -81.16113, -84.32227, -83.9248, -80.41602, -75.95898, -71.20605, 
    -66.35156, -61.42188,
  -76.31348, -80.46484, -83.29004, -82.94727, -79.76465, -75.50098, 
    -70.85645, -66.06738, -61.17969,
  -75.82617, -79.78027, -82.34863, -82.04199, -79.11914, -75.03516, 
    -70.49512, -65.77539, -60.93164,
  -75.29395, -79.05566, -81.40234, -81.125, -78.42773, -74.52441, -70.09668, 
    -65.45215, -60.65723,
  -74.65527, -78.20996, -80.34766, -80.09375, -77.61914, -73.91211, -69.6123, 
    -65.06055, -60.3252,
  -73.79297, -77.10156, -79.0166, -78.78711, -76.55762, -73.08301, -68.94727, 
    -64.52246, -59.86816,
  -72.42383, -75.40137, -77.05469, -76.84961, -74.92969, -71.76562, 
    -67.87012, -63.65137, -59.12402,
  -69.46191, -71.88965, -73.16406, -72.9834, -71.57617, -68.9082, -65.45312, 
    -61.7041, -57.43652 ;

 longitude =
  169.0723, 175.2617, -156.0635, -57.94629, -38.32422, -33.57617, -31.45605, 
    -31.33105, -30.95117,
  150.168, 143.4307, 114.9785, 10.5498, -9.655273, -15.50781, -18.35449, 
    -20.55176, -21.98242,
  141.21, 129.584, 95.69043, 30.51562, 3.101562, -6.956055, -12.01758, 
    -15.39746, -17.6748,
  135.5586, 121.8145, 89.27637, 38.26758, 10.46973, -1.548828, -7.87793, 
    -12.01172, -14.82324,
  131.3408, 116.5332, 85.87402, 42.58984, 15.58203, 2.491211, -4.688477, 
    -9.381836, -12.59277,
  127.7979, 112.4229, 83.59863, 45.55469, 19.63184, 5.892578, -1.925781, 
    -7.083984, -10.62793,
  124.5156, 108.8584, 81.8291, 47.90137, 23.20312, 9.061523, 0.7197266, 
    -4.860352, -8.712891,
  121.1562, 105.4297, 80.27246, 49.99609, 26.68164, 12.32617, 3.524414, 
    -2.477539, -6.641602,
  117.3428, 101.7773, 78.74609, 52.08301, 30.4248, 16.06641, 6.847656, 
    0.3808594, -4.128906,
  112.46, 97.44238, 77.07617, 54.4043, 34.92773, 20.90918, 11.3418, 4.320312, 
    -0.6074219,
  104.8398, 91.32617, 74.91992, 57.45801, 41.38477, 28.57422, 18.96191, 
    11.20215, 5.745117 ;

 lunar_azimuth_angle =
  289.9531, 281.375, 250.0625, 149.0391, 126.25, 118.0703, 112.2344, 
    108.1484, 103.5625,
  307.6328, 312.1016, 338.0469, 79.72656, 96.95312, 99.58594, 98.97656, 
    97.49219, 95.04688,
  316.0312, 325.4453, 356.9062, 59.41406, 83.9375, 90.88281, 92.60938, 
    92.44531, 91,
  321.3203, 332.8984, 3.046875, 51.44531, 76.41406, 85.39062, 88.46875, 
    89.14844, 88.33594,
  325.2578, 337.9297, 6.242188, 46.96094, 71.19531, 81.29688, 85.28125, 
    86.59375, 86.25781,
  328.5625, 341.8281, 8.34375, 43.85938, 67.05469, 77.85156, 82.53906, 
    84.375, 84.4375,
  331.6094, 345.1953, 9.945312, 41.39062, 63.39844, 74.64844, 79.91406, 
    82.23438, 82.67188,
  334.7188, 348.4062, 11.32812, 39.16406, 59.83594, 71.35938, 77.14062, 
    79.94531, 80.77344,
  338.2344, 351.8047, 12.64844, 36.92188, 56, 67.59375, 73.86719, 77.21875, 
    78.47656,
  342.7109, 355.7891, 14.03906, 34.39844, 51.39062, 62.73438, 69.46875, 
    73.48438, 75.28906,
  349.6094, 1.304688, 15.73438, 31.03906, 44.79688, 55.11719, 62.10156, 
    67.05469, 69.625 ;

 lunar_zenith_angle =
  115.9141, 118.2734, 120.4844, 122.5547, 124.5078, 126.2969, 127.7812, 
    129.3359, 130.3984,
  112.4297, 114.7188, 116.8828, 118.8984, 120.7656, 122.4688, 123.9297, 
    125.2891, 126.3047,
  110.6797, 112.9375, 115.0781, 117.0625, 118.8984, 120.5703, 122.0078, 
    123.3047, 124.3047,
  109.4766, 111.7188, 113.8359, 115.8047, 117.625, 119.2734, 120.7031, 
    121.9766, 122.9531,
  108.5156, 110.7422, 112.8438, 114.8047, 116.6094, 118.2422, 119.6562, 
    120.9141, 121.8828,
  107.6406, 109.8594, 111.9531, 113.8984, 115.6953, 117.3125, 118.7188, 
    119.9609, 120.9219,
  106.7812, 108.9844, 111.0625, 112.9922, 114.7812, 116.3906, 117.7891, 
    119.0234, 119.9688,
  105.8203, 108.0156, 110.0781, 111.9922, 113.7656, 115.3672, 116.75, 
    117.9844, 118.9219,
  104.625, 106.7969, 108.8438, 110.7344, 112.5, 114.0938, 115.4531, 116.6953, 
    117.6172,
  102.8672, 105, 107.0234, 108.8906, 110.6562, 112.2266, 113.5625, 114.8203, 
    115.7266,
  99.41406, 101.4688, 103.4219, 105.2266, 107.0547, 108.5703, 109.8438, 
    111.2188, 112.0547 ;

 noise_diode_counts =
  -192255.5, 7.937811e+10, 4.024952e+10, 1.338743e+11, 9.62642e+10, 
    1.051153e+11, 2.48728e+10, 2.748968e+10, -541572, -389927.8, -357267.9, 
    -451875.7,
  -192455, 7.951131e+10, 4.031503e+10, 1.340114e+11, 9.636364e+10, 
    1.052543e+11, 2.492204e+10, 2.752103e+10, -541962.3, -390597.3, 
    -357059.7, -452165,
  -192556.8, 7.952875e+10, 4.030691e+10, 1.34039e+11, 9.642175e+10, 
    1.052789e+11, 2.489782e+10, 2.753012e+10, -541995.4, -390517.7, 
    -357405.7, -452896.7,
  -192567.2, 7.954548e+10, 4.031101e+10, 1.341124e+11, 9.64358e+10, 
    1.05379e+11, 2.49359e+10, 2.755398e+10, -542123.6, -389925.1, -356806.9, 
    -452140.1,
  -192313.8, 7.977819e+10, 4.04354e+10, 1.345669e+11, 9.674735e+10, 
    1.056344e+11, 2.494573e+10, 2.760563e+10, -540990.2, -389929.5, 
    -356355.5, -451428.3,
  -192336.1, 7.986746e+10, 4.047947e+10, 1.346461e+11, 9.684315e+10, 
    1.056485e+11, 2.500115e+10, 2.764812e+10, -541106, -389861.9, -356464.5, 
    -451283.9,
  -192411.4, 7.989448e+10, 4.048347e+10, 1.346543e+11, 9.674249e+10, 
    1.056623e+11, 2.500555e+10, 2.76274e+10, -540893.8, -389571.6, -356420.2, 
    -451078.5,
  -191843.5, 7.995843e+10, 4.049235e+10, 1.347196e+11, 9.686094e+10, 
    1.057265e+11, 2.501101e+10, 2.764078e+10, -539979.1, -389207, -355907.8, 
    -450638.4,
  -191027.5, 8.01557e+10, 4.057723e+10, 1.349386e+11, 9.701532e+10, 
    1.058361e+11, 2.50446e+10, 2.767011e+10, -539616.1, -389281.2, -355800.9, 
    -449215.4 ;

 scAltitude = 513.2554, 514.1388, 514.68, 514.8704, 514.703, 514.2038, 
    513.3773, 512.2527, 510.8646 ;

 scLatitude = -75.80539, -79.76538, -82.34402, -82.06026, -79.13639, 
    -75.04731, -70.51117, -65.77578, -60.93563 ;

 scLongitude = 127.9064, 112.5719, 83.7981, 45.69278, 19.7016, 5.9615, 
    -1.902194, -6.965672, -10.54837 ;

 scPosECEF =
  -1041.255, 1337.243, -6659.007,
  -471.477, 1134.216, -6760.899,
  99.50891, 915.7113, -6809.802,
  667.1064, 683.437, -6805.346,
  1226.729, 439.2711, -6747.562,
  1773.891, 185.2384, -6636.923,
  2304.256, -76.52837, -6474.27,
  2813.58, -343.7532, -6260.881,
  3297.886, -614.1072, -5998.395 ;

 scQuatECEF =
  0.979834, 0.002474682, -0.1079128, 0.1681489,
  0.9817724, 0.01047037, -0.06512038, 0.1782492,
  0.9817343, 0.01868469, -0.02224391, 0.188026,
  0.9797305, 0.0270858, 0.02061385, 0.1974072,
  0.9757617, 0.03570591, 0.06338427, 0.2063897,
  0.9698361, 0.04447604, 0.1060005, 0.2149508,
  0.9619745, 0.05343207, 0.1483336, 0.2230408,
  0.9521869, 0.06252164, 0.1903324, 0.2306613,
  0.9404965, 0.07173561, 0.2319157, 0.2377717 ;

 scRollAngle = 9.988458, 9.997854, 9.993788, 10.00702, 10.01405, 10.01326, 
    10.01118, 10.01077, 10.01045 ;

 scVelECEF =
  7.095409, -2.434456, -1.60188,
  7.139412, -2.637982, -0.9437096,
  7.125648, -2.821125, -0.2781661,
  7.054487, -2.981793, 0.3894352,
  6.926689, -3.118118, 1.053982,
  6.743517, -3.228327, 1.710317,
  6.50671, -3.311056, 2.353408,
  6.218444, -3.364925, 2.978187,
  5.881242, -3.388901, 3.579775 ;

 sensor_azimuth_angle =
  261.6641, 254.3838, 224.6152, 125.4082, 104.6895, 98.83398, 95.61523, 
    94.32031, 92.80469,
  280.2676, 286.0781, 313.5996, 57.10547, 76.38184, 81.29785, 83.21582, 
    84.44922, 84.92969,
  289.1953, 299.9668, 333.0029, 37.3291, 63.8877, 73.08301, 77.29297, 
    79.79395, 81.20605,
  295.0391, 307.9639, 339.6748, 29.87012, 56.8457, 68.03418, 73.55078, 
    76.84473, 78.83887,
  300.1162, 314.0762, 343.8721, 26.3252, 52.47656, 64.70215, 71.06055, 
    74.87891, 77.2793,
  52.11133, 60.99414, 81.15527, 133.3174, 143.3379, 124.8086, 153.2354, 
    90.63184, 95.83691,
  123.0303, 138.1934, 164.7432, 198.2041, 222.415, 236.0586, 243.9111, 
    248.917, 252.2451,
  127.2197, 142.4375, 167.0908, 196.8682, 219.6758, 233.5186, 241.8086, 
    247.2607, 250.8896,
  131.2246, 146.3184, 168.8789, 195.0752, 216.2598, 230.1416, 238.8857, 
    244.8447, 248.8623,
  136.0791, 150.6973, 170.667, 192.9443, 212.0195, 225.6367, 234.8047, 
    241.3906, 245.9072,
  143.4053, 156.6807, 172.8535, 190.085, 205.915, 218.4873, 227.8691, 
    235.332, 240.5518 ;

 sensor_view_angle =
  60.15625, 60.21289, 60.2334, 60.22656, 60.3125, 60.43359, 60.375, 60.86719, 
    60.90039,
  48.09277, 48.15918, 48.1875, 48.15527, 48.23242, 48.37305, 48.30859, 
    48.80469, 48.83105,
  36.04199, 36.09082, 36.13574, 36.07617, 36.14746, 36.29297, 36.22949, 
    36.7373, 36.74023,
  23.98145, 24.01172, 24.07031, 23.99219, 24.06543, 24.20605, 24.14062, 
    24.66699, 24.63281,
  11.90332, 11.93555, 11.99707, 11.91602, 12.00098, 12.13574, 12.05762, 
    12.60352, 12.52441,
  -0.4189453, -0.3759766, -0.3349609, -0.3251953, -0.2744141, 0.2685547, 
    0.2177734, 0.6035156, 0.4833984,
  -12.11328, -12.04492, -11.99805, -12.08691, -12.00977, -11.83398, 
    -11.95801, -11.40527, -11.55859,
  -24.04199, -23.9873, -23.9541, -24.05176, -23.96973, -23.77539, -23.91992, 
    -23.37402, -23.54688,
  -35.99805, -35.99805, -35.98242, -36.07617, -35.9375, -35.77051, -35.91992, 
    -35.37988, -35.55664,
  -47.95312, -48.01367, -48.02148, -48.10059, -47.87695, -47.77832, 
    -47.91504, -47.38867, -47.55859,
  -59.87793, -59.96875, -60.00391, -60.06348, -59.75684, -59.75098, -59.8584, 
    -59.35645, -59.51953 ;

 sensor_zenith_angle =
  69.54883, 69.65332, 69.69629, 69.69141, 69.82031, 69.99902, 69.89062, 
    70.63965, 70.66211,
  53.50684, 53.59668, 53.63672, 53.60059, 53.69238, 53.8584, 53.77148, 
    54.36426, 54.38086,
  39.46289, 39.52441, 39.57812, 39.5127, 39.5918, 39.75391, 39.67676, 
    40.24512, 40.23926,
  26.04297, 26.0791, 26.14648, 26.06152, 26.1416, 26.29395, 26.21875, 
    26.79395, 26.75,
  12.87402, 12.91113, 12.97852, 12.89062, 12.98242, 13.12793, 13.04102, 
    13.63086, 13.54395,
  0.4521484, 0.40625, 0.3613281, 0.3515625, 0.296875, 0.2900391, 0.2353516, 
    0.6523438, 0.5224609,
  13.10156, 13.0293, 12.97949, 13.0752, 12.99219, 12.80078, 12.93457, 
    12.33301, 12.49707,
  26.11035, 26.05371, 26.01855, 26.12695, 26.03613, 25.82031, 25.97656, 
    25.37305, 25.55762,
  39.41309, 39.41992, 39.4043, 39.5127, 39.35449, 39.16309, 39.32715, 
    38.70996, 38.90039,
  53.33887, 53.4209, 53.43652, 53.53418, 53.2627, 53.1377, 53.2959, 52.64746, 
    52.83887,
  69.12598, 69.28223, 69.34766, 69.44434, 68.97266, 68.95508, 69.10156, 
    68.32422, 68.54004 ;

 solar_azimuth_angle =
  7.390625, 0.7890625, 331.8203, 233.5312, 213.8828, 209.2656, 207.4297, 
    207.8516, 208.2109,
  26.44531, 32.625, 60.63281, 164.7578, 184.7891, 190.6172, 193.6016, 
    196.1641, 198.1562,
  35.45312, 46.4375, 79.82031, 144.6172, 171.7812, 181.7422, 186.8594, 
    190.5078, 193.2578,
  41.125, 54.17969, 86.15625, 136.7344, 164.2344, 176.0938, 182.4297, 
    186.7656, 189.9844,
  45.35156, 59.42969, 89.49219, 132.2969, 158.9688, 171.8594, 178.9922, 
    183.8359, 187.3984,
  48.89844, 63.50781, 91.69531, 129.2266, 154.7734, 168.2734, 176.0078, 
    181.2656, 185.1094,
  52.17969, 67.03125, 93.39062, 126.7734, 151.0547, 164.9219, 173.1328, 
    178.7656, 182.8672,
  55.52344, 70.41406, 94.85938, 124.5469, 147.4062, 161.4375, 170.0625, 
    176.0703, 180.4219,
  59.32031, 74, 96.27344, 122.2969, 143.4453, 157.4219, 166.3984, 172.8125, 
    177.4297,
  64.15625, 78.21875, 97.75, 119.7109, 138.6016, 152.1562, 161.3906, 
    168.2578, 173.1797,
  71.63281, 84.04688, 99.47656, 116.0703, 131.4297, 143.6016, 152.6797, 
    160.1328, 165.3203 ;

 solar_beta_angle = 16.36152, 16.6794, 17.00591, 17.33092, 17.64458, 
    17.93662, 18.19846, 18.42097, 18.59702 ;

 solar_zenith_angle =
  80.92969, 85.6875, 90.4375, 95.16406, 99.85156, 104.5, 109.1484, 113.6328, 
    118.1641,
  82.04688, 86.84375, 91.63281, 96.41406, 101.1719, 105.8984, 110.625, 
    115.2656, 119.9062,
  82.61719, 87.42969, 92.23438, 97.03125, 101.8125, 106.5703, 111.3203, 
    116.0234, 120.7109,
  83.01562, 87.82812, 92.64062, 97.44531, 102.2422, 107.0156, 111.7812, 
    116.5078, 121.2266,
  83.34375, 88.15625, 92.96875, 97.78125, 102.5781, 107.3672, 112.1484, 
    116.8906, 121.6328,
  83.63281, 88.44531, 93.26562, 98.07812, 102.8828, 107.6797, 112.4688, 
    117.2266, 121.9766,
  83.92969, 88.74219, 93.55469, 98.36719, 103.1797, 107.9766, 112.7812, 
    117.5469, 122.3203,
  84.25, 89.0625, 93.875, 98.69531, 103.5078, 108.3125, 113.1172, 117.8984, 
    122.6797,
  84.66406, 89.46875, 94.27344, 99.09375, 103.9062, 108.7109, 113.5312, 
    118.3125, 123.1094,
  85.26562, 90.0625, 94.85938, 99.67188, 104.4688, 109.2812, 114.1016, 
    118.8906, 123.7109,
  86.46094, 91.21875, 95.99219, 100.7812, 105.5234, 110.3281, 115.1484, 
    119.8984, 124.7422 ;
}
