netcdf tms_rad_2 {
dimensions:
	spots = 11 ;
	scans = 11 ;
	channels = 12 ;
	cal_spots = 10 ;
	sensors = 6 ;
	coord = 3 ;
	coord2 = 4 ;
variables:
	float AttitudeErrorDeg(spots, scans) ;
		AttitudeErrorDeg:_FillValue = -999.f ;
		AttitudeErrorDeg:long_name = "Estimated Attitude Error" ;
		AttitudeErrorDeg:Description = "Estimated star tracker attitude error magnitude" ;
		AttitudeErrorDeg:units = "deg" ;
		AttitudeErrorDeg:Valid\ Range = 0.f, 180.f ;
	ubyte Day(scans) ;
		Day:_FillValue = 255UB ;
		Day:long_name = "UTC day" ;
		Day:Description = "UTC day of month for the nadir ADC spot." ;
		Day:units = "days" ;
		Day:Valid\ Range = 1UB, 31UB ;
	ubyte Hour(scans) ;
		Hour:_FillValue = 255UB ;
		Hour:long_name = "UTC hour" ;
		Hour:Description = "UTC hour of day for the nadir ADC spot." ;
		Hour:units = "months" ;
		Hour:Valid\ Range = 0UB, 23UB ;
	ushort Millisecond(scans) ;
		Millisecond:_FillValue = 65535US ;
		Millisecond:long_name = "UTC millisecond" ;
		Millisecond:Description = "UTC millisecond of second for the nadir ADC spot." ;
		Millisecond:units = "milliseconds" ;
		Millisecond:Valid\ Range = 0US, 999US ;
	ubyte Minute(scans) ;
		Minute:_FillValue = 255UB ;
		Minute:long_name = "UTC minute" ;
		Minute:Description = "UTC minute of our for the nadir spot." ;
		Minute:units = "minutes" ;
		Minute:Valid\ Range = 0UB, 59UB ;
	ubyte Month(scans) ;
		Month:_FillValue = 255UB ;
		Month:long_name = "UTC month" ;
		Month:Description = "UTC month of year for the nadir ADC spot." ;
		Month:units = "months" ;
		Month:Valid\ Range = 1UB, 12UB ;
	float NEDT_DS(scans, channels) ;
		NEDT_DS:_FillValue = -999.f ;
		NEDT_DS:long_name = "NEDT of cold cal. measurement" ;
		NEDT_DS:units = "K" ;
		NEDT_DS:Valid\ Range = 0.f, 100.f ;
		NEDT_DS:Description = "Estimated  NEDT  using ten samples of deep space.  Used the product of gain  (K/DN),  sample standard deviation  (DN), and normal distribution bias correction (N=10)" ;
	float NEDT_ICT(scans, channels) ;
		NEDT_ICT:_FillValue = -999.f ;
		NEDT_ICT:long_name = "NEDT of internal cal target measurement" ;
		NEDT_ICT:Description = "Estimated NEDT using ten samples viewing the internal calibration target. Used the product of gain (K/DN), sample standard deviation (DN), and normal distribution bias correction (N=10)" ;
		NEDT_ICT:units = "K" ;
		NEDT_ICT:Valid\ Range = 0.f, 100.f ;
	float NEDT_ND(scans, channels) ;
		NEDT_ND:_FillValue = -999.f ;
		NEDT_ND:long_name = "NEDT of hot cal. measurement" ;
		NEDT_ND:Description = "Estimated NEDT using ten samples with noise diode turned on viewing deep space. Used the product of gain (K/DN), sample standard deviation (DN), and normal distribution bias correction (N=10)" ;
		NEDT_ND:units = "K" ;
		NEDT_ND:Valid\ Range = 0.f, 100.f ;
	ubyte NumGPSSats(spots, scans) ;
		NumGPSSats:_FillValue = 255UB ;
		NumGPSSats:long_name = "Number of GPS satellites" ;
		NumGPSSats:Description = "Number of GPS satellites utilized for position calculation." ;
		NumGPSSats:units = "unitless" ;
		NumGPSSats:Valid\ Range = 0UB, 99UB ;
	ubyte Second(scans) ;
		Second:_FillValue = 255UB ;
		Second:long_name = "UTC second" ;
		Second:Description = "UTC second of minute for the nadir ADC spot." ;
		Second:units = "seconds" ;
		Second:Valid\ Range = 0UB, 60UB ;
	ubyte StarTrackerStatus(spots, scans) ;
		StarTrackerStatus:_FillValue = 255UB ;
		StarTrackerStatus:long_name = "Star Tracker Attitude Status Flag" ;
		StarTrackerStatus:Description = "Star Tracker Attitude Status (0=OK,1=Pending,2=Bad,3=Too_Few_Stars)" ;
		StarTrackerStatus:units = "unitless" ;
		StarTrackerStatus:Valid\ Range = 0UB, 25UB ;
	float Ta_ICT(scans, channels) ;
		Ta_ICT:_FillValue = -999.f ;
		Ta_ICT:long_name = "antenna temperature of internal cal target" ;
		Ta_ICT:units = "K" ;
		Ta_ICT:Valid\ Range = 0.f, 400.f ;
		Ta_ICT:Description = "Measured antenna temperature of the internal  calibration target, using the  noise diode as warm  cal source." ;
	ushort Year(scans) ;
		Year:_FillValue = 65535US ;
		Year:long_name = "UTC year" ;
		Year:Description = "UTC year of the nadir ADC spot." ;
		Year:units = "years" ;
		Year:Valid\ Range = 2020US, 2035US ;
	float brightness_temperature(spots, scans, channels) ;
		brightness_temperature:_FillValue = -999.f ;
		brightness_temperature:least_significant_digit = 2LL ;
		brightness_temperature:long_name = "Earth radiometric brightness temperature" ;
		brightness_temperature:units = "K" ;
		brightness_temperature:Valid\ Range = 0.f, 350.f ;
		brightness_temperature:Description = "Planck blackbody equivalent brightness temperatures  resampled to the channel 10  (G3)  boresight-Earth ellipsoid intersection." ;
	float clear_fraction(spots, scans, channels) ;
		clear_fraction:_FillValue = -999.f ;
		clear_fraction:least_significant_digit = 3LL ;
		clear_fraction:long_name = "Clear Fraction" ;
		clear_fraction:units = "Unitless" ;
		clear_fraction:Valid\ Range = 0.f, 1.f ;
		clear_fraction:Description = "Cloud-clear  fraction of each spot from time-matched geostationary satellite cloud mask, weighted by each channel\'s  antenna pattern and resampled to the channel 10  (G3) boresight-Earth ellipsoid intersection." ;
	float cold_target_counts(scans, channels) ;
		cold_target_counts:_FillValue = 0.f ;
		cold_target_counts:long_name = "Cold target counts" ;
		cold_target_counts:Description = "Mean counts (digital number) of the cold (deep space) calibration sector" ;
	ushort combinedQualityFlag(spots, scans, channels) ;
		combinedQualityFlag:_FillValue = 65535US ;
		combinedQualityFlag:long_name = "Combined Quality Flag" ;
		combinedQualityFlag:Description = "Bit 1: reserved, Bit2: non-ocean, Bit 3: Outlier timestamp, Bit 4: RFI, Bit 5: ICT-ND consistency, Bit 6: Attitude Quality, Bit 7: flagICTCal, Bit 8: flagNDCal, Bit 9: flagColdCal, Bit 10: flagPLOrientation, Bit 11: flagDayNight, Bit 12: flagAscDesc, Bit 13: flagManeuver, Bit 14: flagSolarIntrusion, Bit 15: flagLunarIntrusion" ;
		combinedQualityFlag:units = "unitless" ;
		combinedQualityFlag:Valid\ Range = 0US, 65534US ;
	float elevation(spots, scans, channels) ;
		elevation:_FillValue = -9999.f ;
		elevation:least_significant_digit = 1LL ;
		elevation:long_name = "Surface elevation" ;
		elevation:Description = "Surface elevation weighted by each channel\'s antenna pattern" ;
		elevation:units = "m" ;
		elevation:Valid\ Range = -1000.f, 10000.f ;
	ubyte flagAscDesc(spots, scans, channels) ;
		flagAscDesc:_FillValue = 255UB ;
		flagAscDesc:long_name = "Ascending/Descending flag" ;
		flagAscDesc:Description = "1 if in descending portion of orbit, 0 if in ascending portion of orbit." ;
		flagAscDesc:units = "unitless" ;
		flagAscDesc:Valid\ Range = 0UB, 1UB ;
	ubyte flagColdCal(cal_spots, scans, channels) ;
		flagColdCal:_FillValue = 255UB ;
		flagColdCal:long_name = "Cold Calibration Spot Flag" ;
		flagColdCal:Description = "Outlier detection flag for deep space calibration spots." ;
		flagColdCal:units = "unitless" ;
		flagColdCal:Valid\ Range = 0UB, 1UB ;
	ubyte flagDayNight(spots, scans, channels) ;
		flagDayNight:_FillValue = 255UB ;
		flagDayNight:long_name = "Day/Night flag" ;
		flagDayNight:Description = "1 if earth is between the sun and spacecraft, 0 if spacecraft is illuminated by sun." ;
		flagDayNight:units = "unitless" ;
		flagDayNight:Valid\ Range = 0UB, 1UB ;
	ubyte flagICTCal(cal_spots, scans, channels) ;
		flagICTCal:_FillValue = 255UB ;
		flagICTCal:long_name = "Internal Calibration Target Spot Flag" ;
		flagICTCal:Description = "Outlier detection flag for internal calibration target spots." ;
		flagICTCal:units = "unitless" ;
		flagICTCal:Valid\ Range = 0UB, 1UB ;
	ubyte flagICT_ND_Consistency(spots, scans, channels) ;
		flagICT_ND_Consistency:_FillValue = 255UB ;
		flagICT_ND_Consistency:long_name = "Internal Cal Target - Noise Diode Consistency Flag" ;
		flagICT_ND_Consistency:Description = "0 = ICT and ND are consistent, 1 = ND inconsistent with ICT thermistor, 2 = antenna_temperature_ND inconsistent with antenna_temperature_ICT, 3=Both conditions true" ;
		flagICT_ND_Consistency:units = "unitless" ;
		flagICT_ND_Consistency:Valid\ Range = 0UB, 3UB ;
	ubyte flagLunarIntrusion(spots, scans, channels) ;
		flagLunarIntrusion:_FillValue = 255UB ;
		flagLunarIntrusion:long_name = "Lunar intrusion flag" ;
		flagLunarIntrusion:Description = "1 if there is a lunar intrusion into the cold space or noise diode calibration sectors, 0 indicates no intrusion." ;
		flagLunarIntrusion:units = "unitless" ;
		flagLunarIntrusion:Valid\ Range = 0UB, 1UB ;
	ubyte flagManeuver(spots, scans, channels) ;
		flagManeuver:_FillValue = 255UB ;
		flagManeuver:long_name = "Spacecraft maneuver flag" ;
		flagManeuver:units = "unitless" ;
		flagManeuver:Valid\ Range = 0UB, 1UB ;
		flagManeuver:Description = "True if the spacecraft is in an  active  maneuver." ;
	ubyte flagNDCal(cal_spots, scans, channels) ;
		flagNDCal:_FillValue = 255UB ;
		flagNDCal:long_name = "Noise Diode Calibration Spot Flag" ;
		flagNDCal:Description = "Outlier detection flag for noise diode calibration spots." ;
		flagNDCal:units = "unitless" ;
		flagNDCal:Valid\ Range = 0UB, 1UB ;
	ubyte flagNonOcean(spots, scans, channels) ;
		flagNonOcean:_FillValue = 255UB ;
		flagNonOcean:long_name = "Non-ocean Flag" ;
		flagNonOcean:Description = "0 is ocean, 1 is land, coastline, or undefined" ;
		flagNonOcean:units = "unitless" ;
		flagNonOcean:Valid\ Range = 0UB, 1UB ;
	ubyte flagOutlierTimestamp(spots, scans) ;
		flagOutlierTimestamp:_FillValue = 255UB ;
		flagOutlierTimestamp:long_name = "Outlier Timestamp flag" ;
		flagOutlierTimestamp:Description = "1 if original spot time stamp was NaN or deviates more than 10% from expected value. These timestamps are replaced with interpolated values." ;
		flagOutlierTimestamp:units = "unitless" ;
		flagOutlierTimestamp:Valid\ Range = 0UB, 1UB ;
	ubyte flagPLOrientation(spots, scans, channels) ;
		flagPLOrientation:_FillValue = 255UB ;
		flagPLOrientation:long_name = "Payload Orientation flag" ;
		flagPLOrientation:Description = "0 if spacecraft is flying payload-first, 1 if spacecraft flying payload-aft." ;
		flagPLOrientation:units = "unitless" ;
		flagPLOrientation:Valid\ Range = 0UB, 1UB ;
	ubyte flagRFI(spots, scans, channels) ;
		flagRFI:_FillValue = 255UB ;
		flagRFI:long_name = "Radio Frequency Interference Flag" ;
		flagRFI:Description = "1 when either spacecraft or ground-source RFI is detected." ;
		flagRFI:units = "unitless" ;
		flagRFI:Valid\ Range = 0UB, 1UB ;
	ubyte flagSDRTX(spots, scans) ;
		flagSDRTX:_FillValue = 255UB ;
		flagSDRTX:long_name = "Software-defined Radio Transmit Flag" ;
		flagSDRTX:Description = "1 when the software-defined radio on the TMS bus is in transmit mode." ;
		flagSDRTX:units = "unitless" ;
		flagSDRTX:Valid\ Range = 0UB, 1UB ;
	ubyte flagSolarIntrusion(spots, scans, channels) ;
		flagSolarIntrusion:_FillValue = 255UB ;
		flagSolarIntrusion:long_name = "Solar intrusion flag" ;
		flagSolarIntrusion:Description = "1 if there is a solar intrusion into the cold space or noise diode calibration sectors, 0 indicates no intrusion." ;
		flagSolarIntrusion:units = "unitless" ;
		flagSolarIntrusion:Valid\ Range = 0UB, 1UB ;
	float instrTemp(sensors, scans) ;
		instrTemp:_FillValue = -999.f ;
		instrTemp:long_name = "Average instrument temperature" ;
		instrTemp:units = "degree Celsius" ;
		instrTemp:Valid\ Range = -50.f, 50.f ;
		instrTemp:Description = "1st:  The W/F RFE temperature; 2nd:  The G-band RFE temperature, 3-6:  ICT  thermistor temperatures." ;
	float internal_cal_target_counts(scans, channels) ;
		internal_cal_target_counts:_FillValue = 0.f ;
		internal_cal_target_counts:long_name = "Internal Calibration Target counts" ;
		internal_cal_target_counts:Description = "Mean counts (digital number) of the internal calibration target sector" ;
	float land_fraction(spots, scans, channels) ;
		land_fraction:_FillValue = -999.f ;
		land_fraction:least_significant_digit = 3LL ;
		land_fraction:long_name = "Land Fraction" ;
		land_fraction:units = "Unitless" ;
		land_fraction:Valid\ Range = 0.f, 1.f ;
		land_fraction:Description = "Land fraction weighted by each  channel\'s antenna pattern, resampled to the channel  10  (G3) boresight-Earth ellipsoid intersection." ;
	float latitude(spots, scans) ;
		latitude:_FillValue = -999.f ;
		latitude:least_significant_digit = 3LL ;
		latitude:long_name = "Latitude: line-of-sight to Earth intersection" ;
		latitude:Description = "Geodetic latitude of the line-of-sight intersection point with the Earth for each spot. Negative values are South. These correspond to the middle of each spots integration period. WGS84" ;
		latitude:units = "degree_north" ;
		latitude:Valid\ Range = -90.f, 90.f ;
	float longitude(spots, scans) ;
		longitude:_FillValue = -999.f ;
		longitude:least_significant_digit = 3LL ;
		longitude:long_name = "Longitude: line-of-sight to Earth intersection" ;
		longitude:Description = "Geodetic longitude of the line-of-sight intersection point with the Earth for each spot. Negative values are West. These correspond to the middle of each spots integration period. WGS84" ;
		longitude:units = "degree_east" ;
		longitude:Valid\ Range = -180.f, 180.f ;
	float lunar_azimuth_angle(spots, scans) ;
		lunar_azimuth_angle:_FillValue = -999.f ;
		lunar_azimuth_angle:long_name = "Line-of-sight lunar azimuth angle" ;
		lunar_azimuth_angle:Description = "The angle between the local north vector at the LOS\'s earth intersection point and a vector pointing at the center of the Moon." ;
		lunar_azimuth_angle:units = "degree" ;
		lunar_azimuth_angle:Valid\ Range = 0.f, 360.f ;
	float lunar_zenith_angle(spots, scans) ;
		lunar_zenith_angle:_FillValue = -999.f ;
		lunar_zenith_angle:long_name = "Line-of-sight lunar zenith angle" ;
		lunar_zenith_angle:Description = "The angle between the local zenith at the LOS\'s earth intersection point and a vector pointing at the center of the Moon." ;
		lunar_zenith_angle:units = "degree" ;
		lunar_zenith_angle:Valid\ Range = 0.f, 180.f ;
	float noise_diode_counts(scans, channels) ;
		noise_diode_counts:_FillValue = 0.f ;
		noise_diode_counts:long_name = "Noise diode counts" ;
		noise_diode_counts:Description = "Mean counts (digital number) of the noise diode calibration sector" ;
	float scAltitude(scans) ;
		scAltitude:_FillValue = -99999.f ;
		scAltitude:long_name = "Spacecraft altitude" ;
		scAltitude:units = "km" ;
		scAltitude:Valid\ Range = 0.f, 1000.f ;
		scAltitude:Description = "The altitude of the spacecraft above the   WGS84  ellipsoid." ;
	float scLatitude(scans) ;
		scLatitude:_FillValue = -999.f ;
		scLatitude:long_name = "Spacecraft latitude" ;
		scLatitude:Description = "The latitude of the spacecraft sub-satellite point. WGS84. " ;
		scLatitude:units = "degrees_north" ;
		scLatitude:Valid\ Range = -90.f, 90.f ;
	float scLongitude(scans) ;
		scLongitude:_FillValue = -999.f ;
		scLongitude:long_name = "Spacecraft longitude" ;
		scLongitude:Description = "The longitude of the spacecraft sub-satellite point. WGS84. " ;
		scLongitude:units = "degrees_east" ;
		scLongitude:Valid\ Range = -180.f, 180.f ;
	float scPosECEF(scans, coord) ;
		scPosECEF:_FillValue = -99999.f ;
		scPosECEF:long_name = "Spacecraft ECEF position" ;
		scPosECEF:Description = "The spacecraft position in ECEF coordinate system.  The first dimension is [x,y,z]. WGS84. Uses 41st ADC spot in each scan for timestamp." ;
		scPosECEF:units = "km" ;
		scPosECEF:Valid\ Range = -10000.f, 10000.f ;
	float scQuatECEF(scans, coord2) ;
		scQuatECEF:_FillValue = -999.f ;
		scQuatECEF:long_name = "Spacecraft Body-to-ECEF quaternion" ;
		scQuatECEF:Description = "The unit length quaternion that rotates from spacecraft body coordinate system to ECEF coordinate system.  The second dimension is [i,j,k,r], where r is the scalar element of the quaternion. WGS84. Uses 41st ADC spot in each scan for timestamp." ;
		scQuatECEF:units = "norm one" ;
		scQuatECEF:Valid\ Range = -1.f, 1.f ;
	float scRollAngle(scans) ;
		scRollAngle:_FillValue = -999.f ;
		scRollAngle:long_name = "Roll angle of the spacecraft" ;
		scRollAngle:Description = "Zero degrees means the spacecraft body Z-axis is aligned with nadir in the spacecraft body XY plane" ;
		scRollAngle:units = "degrees" ;
		scRollAngle:Valid\ Range = 0.f, 360.f ;
	float scVelECEF(scans, coord) ;
		scVelECEF:_FillValue = -99999.f ;
		scVelECEF:long_name = "Spacecraft ECEF velocity" ;
		scVelECEF:Description = "The spacecraft velocity in ECEF coordinate system.  The first dimension is [x,y,z]. WGS84. Uses 41st ADC spot in each scan for timestamp." ;
		scVelECEF:units = "km/s" ;
		scVelECEF:Valid\ Range = -10.f, 10.f ;
	float sensor_azimuth_angle(spots, scans) ;
		sensor_azimuth_angle:_FillValue = -999.f ;
		sensor_azimuth_angle:long_name = "Line-of-sight azimuth angle" ;
		sensor_azimuth_angle:units = "degree" ;
		sensor_azimuth_angle:Valid\ Range = 0.f, 360.f ;
		sensor_azimuth_angle:Description = "The angle between the local north vector at the  LOS earth intersection point and the inverse  LOS vector  (a vector pointing toward the satellite from earth)." ;
	float sensor_view_angle(spots, scans) ;
		sensor_view_angle:_FillValue = -999.f ;
		sensor_view_angle:long_name = "Line-of-sight scan angle" ;
		sensor_view_angle:Description = "The scan angle between the satellite local nadir and the Line-Of-Sight (LOS) vector from radiometer aperture." ;
		sensor_view_angle:units = "degree" ;
		sensor_view_angle:Valid\ Range = -180.f, 180.f ;
	float sensor_zenith_angle(spots, scans) ;
		sensor_zenith_angle:_FillValue = -999.f ;
		sensor_zenith_angle:long_name = "Line-of-sight zenith angle" ;
		sensor_zenith_angle:Description = "The angle between the local zenith at the LOS earth intersection point and the inverse LOS vector (a vector pointing toward the satellite from earth)." ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:Valid\ Range = 0.f, 90.f ;
	float solar_azimuth_angle(spots, scans) ;
		solar_azimuth_angle:_FillValue = -999.f ;
		solar_azimuth_angle:long_name = "Line-of-sight solar azimuth angle" ;
		solar_azimuth_angle:Description = "The angle between the local north vector at the LOS\'s earth intersection point and a vector pointing at the center of the Sun." ;
		solar_azimuth_angle:units = "degree" ;
		solar_azimuth_angle:Valid\ Range = 0.f, 360.f ;
	float solar_beta_angle(scans) ;
		solar_beta_angle:_FillValue = -999.f ;
		solar_beta_angle:long_name = "Solar beta angle" ;
		solar_beta_angle:units = "degree" ;
		solar_beta_angle:Valid\ Range = -90.f, 90.f ;
		solar_beta_angle:Description = "The angle the satellite-sun  vector extends out of the orbital plane. Uses  41st  ADC  spot in each scan for timestamp." ;
	float solar_zenith_angle(spots, scans) ;
		solar_zenith_angle:_FillValue = -999.f ;
		solar_zenith_angle:long_name = "Line-of-sight solar zenith angle" ;
		solar_zenith_angle:Description = "The angle between the local zenith at the LOS\'s earth intersection point and a vector pointing at the center of the Sun." ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:Valid\ Range = 0.f, 180.f ;

// global attributes:
		:processing_stream = "NRT" ;
		:SV_ID = 2LL ;
		:PL_ID = 3LL ;
		:DataSetQuality = "Validated" ;
		:satellite_sub_identifier = 102LL ;
		:L1BR_SW_Ver = "1.0" ;
		:version = "V01-00" ;
		:CloudMaskFiles = "MSG3-SEVI-MSGCLMK-0100-0100-20250915003000.000000000Z-NA" ;
		:Filename = "TMS02.1B-TBR.V01-00.NRT.ST20250915-002225.ET20250915-003601.CT20250915-013139.nc" ;
		:L1B_file = "TMS02.1B-TB.V01-00.NRT.ST20250915-002225.ET20250915-003601.CT20250915-013123.nc" ;
		:create_time = "2025-09-15T01:31:39" ;
		:start_time = "2025-09-15T00:22:25" ;
		:end_time = "2025-09-15T00:36:01" ;
		:platform = "Tomorrow-S02" ;
		:collection = "TS02_L1B-TBR" ;
		:history = "Wed Jan 14 20:06:24 2026: ncks -d scans,0,,40 -d spots,0,,8 /home/Yaping.Wang/scratchda/TMS/TS02_L1B-TBR/20250915/TMS02.1B-TBR.V01-00.NRT.ST20250915-002225.ET20250915-003601.CT20250915-013139.nc tms_rad_2_thin.nc" ;
		:NCO = "netCDF Operators version 5.2.4 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 AttitudeErrorDeg =
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537,
  0.1495085, 0.01164382, 0.01118997, 0.01139705, 0.01726123, 0.01121239, 
    0.01104035, 0.009431244, 0.007883956, 0.006455775, 0.009790537 ;

 Day = 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15 ;

 Hour = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Millisecond = 550, 542, 544, 543, 543, 544, 544, 544, 544, 547, 545 ;

 Minute = 22, 23, 25, 26, 27, 29, 30, 31, 33, 34, 35 ;

 Month = 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9 ;

 NEDT_DS =
  1.001624, 0.5173188, 0.5526987, 0.3812869, 0.2667916, 0.2818989, 0.63255, 
    0.6099188, 0.4337778, 0.5121636, 0.295386, 0.2189684,
  0.5619661, 0.3528214, 0.4848758, 0.2560758, 0.4909678, 0.2931798, 
    0.5144768, 0.438102, 0.3091479, 0.5638668, 0.3073961, 0.5316757,
  0.8754088, 0.3050126, 0.5748503, 0.2409612, 0.3417832, 0.2759507, 
    0.5181042, 0.623458, 0.4719745, 0.1822471, 0.2522821, 0.3648341,
  0.724678, 0.2649715, 0.3850203, 0.3684633, 0.407885, 0.3369833, 0.4385249, 
    0.6761729, 0.537834, 0.5362627, 0.1952811, 0.5026918,
  1.092921, 0.351221, 0.407772, 0.368641, 0.3542533, 0.3947842, 0.5315484, 
    0.4824981, 0.400079, 0.2489985, 0.3758078, 0.5561579,
  0.9997575, 0.3491934, 0.2824631, 0.4293742, 0.3044716, 0.4368702, 
    0.8023921, 0.7320461, 0.2826692, 0.288022, 0.152255, 0.4212469,
  0.9796449, 0.2907054, 0.439433, 0.5340598, 0.3876022, 0.2902304, 0.4512801, 
    0.5803837, 0.3371436, 0.3714224, 0.3628784, 0.4777229,
  1.230549, 0.3607419, 0.3167986, 0.3967812, 0.3200733, 0.4273889, 0.524421, 
    0.6783041, 0.446292, 0.4206127, 0.465693, 0.6216232,
  1.247702, 0.2894045, 0.3041876, 0.3318314, 0.4111099, 0.5101196, 0.4426977, 
    0.7559478, 0.4425943, 0.224205, 0.2978128, 0.4758202,
  1.443404, 0.3046812, 0.3914818, 0.252068, 0.3401738, 0.375342, 0.5546524, 
    0.589788, 0.4202082, 0.6704779, 0.1968301, 0.4504799,
  0.6861798, 0.3955182, 0.368647, 0.3069108, 0.5562314, 0.3696519, 0.5245993, 
    0.3738413, 0.4304441, 0.424659, 0.2453691, 0.4627856 ;

 NEDT_ICT =
  0.6861477, 0.5750291, 0.767269, 0.3895918, 0.4581232, 0.6033235, 1.102908, 
    1.188643, 0.5336213, 0.3448062, 0.4622908, 0.715323,
  1.209891, 0.6057532, 0.8490434, 0.3828416, 0.5823827, 0.7239244, 1.477338, 
    1.469795, 0.5088533, 0.4344633, 0.3472328, 0.5139511,
  1.249888, 0.5408154, 0.6020073, 0.3505194, 0.5127651, 0.5509431, 0.7872076, 
    0.98557, 0.4226561, 0.2967516, 0.4611303, 0.3756003,
  0.9188416, 0.3863249, 0.6800685, 0.4037109, 0.5461495, 1.039775, 1.245417, 
    1.016632, 0.5268353, 0.4013506, 0.3895041, 0.5334399,
  0.6740161, 0.4917101, 0.4435677, 0.3157335, 0.7442091, 0.7243821, 
    0.9479706, 0.815642, 0.561743, 0.2889254, 0.3379302, 0.3346155,
  1.158988, 0.5163754, 0.5612075, 0.5795678, 0.8386697, 0.6991135, 1.089278, 
    0.7599811, 0.454466, 0.481936, 0.4233983, 0.6899376,
  0.7081535, 0.3059663, 0.6530881, 0.6548563, 0.6962439, 0.732612, 1.330453, 
    1.058651, 0.5980603, 0.4039768, 0.3765013, 0.4510728,
  0.6540409, 0.3968158, 0.7275361, 0.6262101, 0.780469, 0.4104654, 0.9845763, 
    1.274026, 0.5584248, 0.5276684, 0.4564299, 1.076677,
  1.157434, 0.4149944, 0.9400972, 0.5214029, 0.7006083, 0.7544192, 0.911677, 
    1.124984, 0.3416553, 0.3733354, 0.5287269, 0.6903161,
  0.8937055, 0.6700594, 0.478474, 0.4141919, 0.7050973, 0.4762555, 0.9407046, 
    0.7797958, 0.4575673, 0.3745311, 0.231132, 0.7179741,
  1.019467, 0.2974453, 0.4049892, 0.6409066, 0.6111615, 0.7981709, 1.257785, 
    0.7790035, 0.5183294, 0.4332817, 0.538719, 1.130336 ;

 NEDT_ND =
  1.34476, 0.6024402, 0.5956612, 0.6036791, 0.7972662, 0.5754913, 0.6934252, 
    0.8911251, 0.6745696, 0.5714796, 0.6196491, 0.6678029,
  0.7750096, 0.4904619, 0.8451681, 0.6702969, 0.7288525, 0.6086602, 
    0.8023472, 0.8122864, 0.90444, 0.7165329, 0.3085068, 0.6127807,
  1.43924, 0.6461712, 0.6832363, 0.558899, 0.6470409, 0.6801497, 1.043007, 
    0.5449768, 0.6461897, 0.3942968, 0.3036317, 0.6076032,
  0.5850706, 0.5038905, 0.4198263, 0.6140941, 0.3829292, 0.7928169, 
    0.5941856, 0.8335512, 0.4858335, 0.4340405, 0.4344335, 0.4955783,
  0.9916829, 0.5048925, 0.3040966, 0.6517109, 0.5936998, 0.4774022, 
    0.8535702, 0.6070156, 0.7580183, 0.4979925, 0.368929, 0.5704895,
  0.9956716, 0.4920812, 0.3631007, 0.5594918, 0.7416469, 0.539224, 0.6152157, 
    0.844448, 0.4691874, 0.6619383, 0.3664509, 0.4919133,
  0.8211234, 0.6422088, 0.6803269, 0.4887806, 0.6043409, 0.6887154, 
    0.8656776, 0.9376606, 0.9392521, 0.8487545, 0.4562739, 0.7729504,
  1.025161, 0.4439862, 0.8150094, 0.5494809, 0.5707206, 0.5673776, 1.200213, 
    0.6527228, 0.4356642, 0.5304946, 0.5556932, 0.6871255,
  0.9868152, 0.4143054, 0.5329369, 0.3434992, 0.477744, 0.5101349, 0.7022565, 
    0.5884613, 0.2462265, 0.4657406, 0.3617439, 0.4811991,
  0.7019104, 0.3691069, 0.6477129, 0.6934158, 0.7809222, 0.6612807, 1.333238, 
    0.7496091, 0.4169885, 0.5040442, 0.395096, 0.9726512,
  0.7216556, 0.8005989, 0.5618867, 0.3613731, 0.6458986, 0.507395, 0.9972363, 
    0.4751005, 0.3231545, 0.4581602, 0.3689879, 0.5083041 ;

 NumGPSSats =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Second = 26, 46, 6, 26, 46, 6, 26, 46, 6, 26, 46 ;

 StarTrackerStatus =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Ta_ICT =
  _, 285.6562, 286.2178, 286.4881, 285.9112, 286.085, 285.805, 286.2158, 
    287.4471, 284.1303, _, 272.1224,
  282.777, 284.3977, 285.2893, 285.0783, 284.944, 285.1229, 284.5701, 
    284.6201, 285.6327, 283.1313, 280.7184, 271.0082,
  282.0461, 284.5019, 285.4126, 284.5728, 285.3122, 284.4119, 284.7183, 
    284.9085, 285.3029, 282.1656, 280.6893, 270.5081,
  282.3474, 284.4267, 285.7307, 284.9407, 285.381, 284.5009, 284.4611, 
    284.3311, 285.1732, 283.3815, 279.7367, 271.4065,
  281.4855, 283.058, 284.0971, 283.78, 284.0175, 283.7225, 283.5349, 283.505, 
    284.9975, 281.1031, 278.9595, 270.2981,
  280.4592, 282.1385, 283.1367, 282.9955, 283.0762, 282.5719, 282.7644, 
    283.2435, 284.0798, 280.7729, 278.5934, 268.549,
  280.1816, 281.5814, 283.3776, 282.5204, 282.268, 282.2647, 282.7281, 
    281.9056, 283.7293, 281.0608, 278.483, 268.7114,
  279.7392, 280.2432, 281.1105, 280.7597, 280.6969, 281.213, 280.8127, 
    281.3635, 282.8283, 279.888, 277.6734, 268.7159,
  279.2215, 280.1213, 281.3953, 280.571, 280.6786, 281.007, 279.8048, 
    280.5279, 282.0269, 278.1347, 276.6116, 266.7681,
  277.1888, 279.8883, 281.3112, 280.705, 280.4748, 280.4326, 279.6497, 
    280.2234, 280.9256, 278.4487, 275.9297, 266.3344,
  276.8598, 279.2366, 280.3836, 279.6516, 279.8475, 279.4813, 279.5412, 
    278.5201, 281.1715, 278.5041, 276.0109, 267.8394 ;

 Year = 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025, 2025 ;

 brightness_temperature =
  204.2812, 241.4531, 238.8125, 229.625, 218.1406, 213.3594, 213.625, 
    224.6016, 239.3672, 254.0156, 262.0625, 265.1719,
  210.6406, 245.8906, 241.2266, 232.9688, 223.6953, 217.3516, 218.6172, 
    224.6484, 248.9141, 259.6797, 264.7578, 267.5391,
  232.0078, 252.3672, 245.3203, 235.2734, 225.9141, 219.8203, 218.6172, 
    225.9375, 252.7656, 261.9141, 268.1641, 271.0781,
  226.7578, 253.625, 246.3047, 237.0078, 225.8359, 218.4062, 217.3125, 
    222.9453, 235.4688, 251.6328, 265.1484, 271.2578,
  225.3359, 256.25, 249.375, 238.3594, 225.5234, 216.7109, 214.0391, 
    221.8984, 228.9609, 246.7422, 263.5156, 274.5547,
  262.0469, 263.3047, 252.5859, 239.8906, 225.3047, 214.3516, 212.2031, 
    221.7344, 232.4453, 255.1797, 267.6719, 274.8047,
  250.8047, 264.0547, 254.0312, 240.1484, 224.4531, 210.9062, 209.6328, 
    221.8594, 239.1484, 263.1562, 274.8125, 280.6406,
  262.9297, 265.5078, 254.5625, 241.4844, 224.7266, 210.6406, 208.6562, 
    221.9531, 243.2109, 265.1094, 277.3516, 281.6641,
  268.7422, 267.9062, 256.4297, 242.5469, 224.4375, 209.5234, 206.2266, 
    221.0391, 243.3672, 263.3594, 273.5312, 282.4375,
  264.0391, 268.1406, 257.5781, 242.7734, 224.75, 209.3125, 206.6406, 
    222.5156, 238.0312, 259.2109, 272.4922, 281.8984,
  274.4062, 270.2812, 258.4688, 243.0781, 223.7344, 210.0156, 205.5781, 
    221.5938, 237.6484, 258.75, 273.7578, 282.0547,
  199.75, 239.0312, 243.5391, 237.5938, 226.3359, 212.8906, 209.0312, 
    219.0078, 243.3594, 256.2109, 263.7031, 264.2969,
  195.8047, 240.2422, 244.4844, 239.6016, 229.0547, 217.5391, 215.2969, 
    221.6406, 248.0156, 259.7031, 267.3438, 266.6719,
  205.9766, 246.0234, 247.5469, 243.0234, 231.0078, 221.6484, 218.1328, 
    223.2109, 258.3516, 266.5156, 271.8828, 272.4375,
  219.0234, 250.9609, 251.1953, 244.4297, 234.0625, 223.6797, 217.4766, 
    222.1875, 256.4609, 262.7656, 267.7734, 271.7109,
  212.8672, 251.3984, 254.0547, 247.6016, 235.3203, 225.7266, 218.4844, 
    222.6797, 236.7734, 250.375, 263.6016, 271.8594,
  228.8906, 258.1016, 257.4453, 249.7578, 235.8203, 220.2344, 214.5859, 
    220.2812, 236.3594, 253.5859, 264.8594, 274.2812,
  240.7266, 265.6719, 262.3125, 253.1484, 236.6953, 220.9219, 209.7891, 
    218.8281, 243.7422, 264.375, 273.5781, 280.5391,
  240.5625, 264.6719, 262.2344, 252.6172, 238.2578, 218.0234, 208.2109, 
    217.7734, 248.5547, 270.1719, 280.3594, 282.125,
  234.7734, 264.3516, 262.5625, 254.6953, 237.3359, 217.3984, 206.4922, 
    217.6172, 249.8516, 269.7656, 280.8359, 287.7109,
  246.4375, 269.3984, 265.9453, 255.2344, 238.6719, 219.7891, 206.5859, 
    216.3281, 244.5703, 265.9453, 278.1562, 286.5391,
  247.625, 270.0938, 265.9297, 255.6484, 238.9531, 217.6953, 206.7656, 
    219.5312, 246.5156, 265.7812, 278.9062, 287.1094,
  208.7109, 240.7969, 244.2344, 241.9609, 229.8438, 216.2344, 208.4922, 
    217.4531, 242.0391, 255.8125, 264.1016, 262.7422,
  216.6562, 244.7578, 248.5547, 244.75, 233.0234, 220.1016, 214.5312, 
    219.7734, 250.0078, 261.3828, 268.0469, 265.8203,
  204.8594, 243.3125, 248.3672, 246.8438, 235.8203, 224.4688, 219.2266, 
    222.2266, 257.8438, 268, 272.2578, 268.0703,
  206.6016, 245.4453, 250.4375, 246.1953, 236.5938, 226.9922, 219.1328, 
    221.8359, 257.4141, 263.8359, 268.0781, 271.9375,
  210.4922, 247.0078, 253.2266, 248.8672, 239.2188, 228.3516, 220.3906, 
    223.8281, 255.5391, 266.0312, 270.7578, 273.2266,
  206.3906, 248.125, 253.2734, 250.8359, 240.8828, 227.0938, 216.0703, 
    218.9531, 243.3594, 253.8281, 265.1172, 274.7031,
  226.7266, 259.7656, 261.1875, 256.6641, 242.8438, 225.3047, 212.8047, 
    217.5156, 248.5156, 264.8516, 273.2969, 281.0312,
  228.1172, 260.5625, 261.8281, 256.8828, 243.6172, 223.6875, 208.4141, 
    217.3984, 252.1328, 271.8125, 280.5, 285.8672,
  232.7266, 264, 265.5391, 259.0547, 244.4453, 224.9609, 209.1172, 215.3828, 
    254.4531, 271.9844, 280.4609, 286.7188,
  242.4766, 266.8828, 268.1797, 260.6406, 245.4062, 223.9688, 209.5078, 
    215.8438, 250.9297, 270.6484, 282.1641, 287.9375,
  241.2578, 268.4922, 267.5625, 261.9688, 244.9766, 224.8828, 208.3125, 
    216.6406, 250.1875, 268.1484, 279.7734, 287.0391,
  213.9922, 241.0781, 245.6094, 244.4688, 233.8984, 216.7656, 209.1875, 214, 
    251.6484, 265.7656, 269.7734, 263.9688,
  212.2344, 241.9219, 248.4531, 245.9844, 236.0938, 222.7812, 213.2734, 
    219.5391, 250.2969, 261.7422, 268.3516, 262.375,
  216.6328, 244.9219, 249.6094, 247.5469, 237.9141, 226.6719, 218.8203, 
    221.5, 254.6953, 264.3984, 270.4766, 266.7188,
  208.5703, 242.5234, 248.6328, 247.375, 239.6953, 228.7188, 220.8281, 
    222.1641, 258.4219, 264.3438, 269.1953, 269.8672,
  213.7266, 245.1719, 250.7812, 250.25, 241.0234, 230.2812, 221.3672, 
    221.2031, 255.9219, 264.8359, 270.2656, 271.1328,
  225.5391, 251.8125, 255.3594, 253.1797, 243.6797, 229, 217.5391, 218.5391, 
    259.9141, 267.4844, 271.6719, 274.5781,
  240.5859, 263.1797, 263.3672, 258.5781, 245.0391, 229.2812, 215.1875, 
    217.8281, 256.0391, 266.5156, 272.3516, 278.0938,
  224.7422, 257.3594, 262.6953, 258.1719, 246.5469, 227.4062, 211.3516, 
    216.2266, 254.9062, 272.2656, 281.5312, 286.1719,
  238.5, 265.5, 266.9922, 261.9297, 247.4062, 227.7266, 210.6562, 215.3125, 
    255.4297, 270.1484, 280.3672, 285.3359,
  243.2266, 267.4375, 266.6328, 261.6328, 248.6719, 227.125, 207.9453, 
    214.8438, 255.5625, 271.9531, 281.4844, 287.4766,
  240.4844, 267.5312, 266.6641, 263.3516, 249.5859, 226.8672, 210.1406, 
    216.8984, 251.4688, 267.7812, 279.5234, 287.2109,
  214.8203, 239.9922, 246.0859, 244.2266, 234.6719, 218.8359, 209.3594, 
    214.5781, 259.2891, 271.4453, 270.5156, 258.8047,
  216.2344, 243.9922, 248.0547, 246.9531, 236.7812, 224.2422, 214.25, 
    219.7344, 249.1328, 260.6016, 268.4219, 263.3047,
  219.3906, 245.0078, 249.3672, 247.5234, 239.1641, 225.6719, 220.4453, 
    222.0781, 252.4922, 261.4609, 269.3828, 264.5391,
  212.0781, 242.2422, 249.0938, 248.8906, 241.2188, 230.1562, 222.4922, 
    220.8438, 257.6016, 262.7969, 268.5625, 267.5938,
  208.4766, 243.0156, 250.1172, 249.3906, 242.4766, 230.9219, 222.2578, 
    221.3203, 255.3594, 265.7812, 270.8672, 268.8438,
  212.8906, 246.8203, 253.0938, 252.4688, 244.0547, 230.4375, 219.5938, 
    220.6094, 261.7812, 269.0312, 273.4297, 274.7969,
  231.4531, 257.9688, 259.9922, 258.8516, 247.875, 229.7578, 215.6094, 
    218.2969, 259.75, 267.9531, 273.0859, 280.5625,
  222.6328, 256.7656, 260.5703, 258.4766, 248.4375, 229.4375, 212.5781, 
    214.9531, 252.875, 270.0078, 280.3359, 284.6328,
  233.9453, 262.7344, 265.9219, 261.3906, 250.3281, 229.9141, 211.6406, 
    215.0938, 253.7891, 270.3281, 279.5547, 285.4062,
  236.6875, 264.8125, 267.2031, 262.6484, 250.9688, 232.1875, 212.9844, 
    215.1094, 256.0078, 273.5781, 282.2969, 288.5156,
  241.8281, 266.3359, 267.6562, 263.6172, 251.2656, 229.6406, 209.4453, 
    215.4844, 252.125, 267.8047, 278.4375, 285.3828,
  211.7812, 240.0781, 246.3984, 245.5078, 235.5938, 219.5703, 206.7969, 
    214.8828, 262.8516, 272.6484, 271.9375, 259.7656,
  218.8281, 244.2266, 247.9062, 246.8594, 236.2578, 221.8828, 212.8359, 
    219.0312, 248.7656, 258.8594, 266.625, 262.4922,
  232.7188, 251.5078, 252.9141, 248.5859, 239.4609, 226.7422, 220.2969, 
    221.75, 253.0078, 262.1094, 270.5, 269.6328,
  215.4219, 244.7734, 249.8828, 248.0156, 240.4219, 230.0234, 223.9219, 
    222.0703, 254.5391, 260.6875, 267.6797, 267.6562,
  205.6719, 239.7188, 247.3047, 248.4375, 242.7344, 231.8828, 221.6953, 
    221.7109, 250.8828, 262.9453, 270.7891, 265.5547,
  214.4766, 246.8516, 253.875, 253.5625, 244.8203, 230.9609, 217.2812, 
    217.4688, 260.9609, 269.2812, 274.5234, 274.2266,
  246.4453, 263.3984, 263.2266, 258.6328, 247.7812, 231.0078, 217.1016, 
    218.1875, 262.3281, 269.6875, 273.875, 278.8281,
  232.3047, 259.4609, 262.7422, 258.9609, 248.8828, 229.3828, 213.2969, 
    216.3984, 254.25, 270.3828, 278.9375, 283.5156,
  228.9062, 260.3828, 263.0859, 262.2812, 250.3125, 230.8906, 213.2266, 
    214.3203, 254.6719, 270.0234, 279.9844, 286.6562,
  234.1562, 262.1484, 264.6484, 263.1328, 251.1094, 230.1406, 213.0938, 
    214.3125, 255.2578, 272.6172, 282.4609, 288.4219,
  238.9766, 265.3906, 267.4297, 263.7422, 251.8516, 230.7578, 211.0625, 
    215.2734, 252.2031, 268.9219, 279.3594, 286.9453,
  208.2109, 238.8516, 246.7812, 246.2578, 234.6484, 218.0703, 207.7656, 
    213.1328, 263.9531, 272.875, 271.9141, 258.125,
  215.0469, 242.3672, 247.6172, 246.2109, 236.6172, 222.0938, 213.1719, 
    216.5703, 248.0391, 258.2656, 266.8672, 262.3203,
  215.8594, 245.0391, 249.5156, 247.6562, 239.6953, 226.3828, 221.3125, 
    221.0156, 253.5, 264.3359, 270.4062, 264.4922,
  215.1875, 244.3594, 248.3672, 247.75, 240.4609, 230.3125, 222.3281, 
    221.7734, 252.5547, 259.5859, 266.7812, 266.7656,
  203.6406, 239.3906, 248.4531, 248.1719, 242.5781, 231.8516, 223.9609, 
    222.0469, 251.3594, 262.9766, 270.7812, 265.2031,
  221.1875, 250, 254.3984, 253.3516, 243.7656, 229.6484, 219.5547, 217.7266, 
    257.6562, 264.8672, 270.7344, 272.5703,
  241.4922, 262, 263.1094, 258.5625, 245.2656, 231.0078, 215.4844, 217.8125, 
    263.4141, 272.7578, 276.0859, 282.4219,
  237.0625, 261.0391, 263.0703, 258.7109, 248.5938, 229.8906, 212.9609, 
    216.4297, 260.875, 273.0859, 279.1172, 283.4922,
  229.7344, 260.8828, 263.25, 261.75, 250.2344, 230.3281, 211.6406, 216.7031, 
    252.9844, 269.9688, 280.1484, 286.6094,
  232.7656, 261.0156, 264.9297, 262.9531, 250.7656, 230.9531, 210.8359, 
    215.1562, 255.9062, 271.5781, 282.0625, 289.0391,
  238.3047, 266.7969, 267.6406, 263.1875, 250.4922, 229.5391, 209.0156, 
    214.6641, 251.3672, 268.5469, 278.7422, 285.6953,
  203.8516, 238.8672, 244.8906, 242.7578, 231.4766, 216.8047, 204.625, 
    213.2656, 261.1094, 271.5156, 271.7969, 260.7578,
  219.9766, 244.5938, 247.7422, 244.875, 234.8281, 220.1641, 212.3438, 
    218.7422, 245.4219, 256.4453, 265.5, 264.1875,
  210.2734, 243.1875, 248.1562, 246.4922, 237.3047, 226.2109, 220.5859, 
    223.0859, 252.3516, 262.2188, 269.1641, 267.2656,
  215.9297, 245.3516, 248.8047, 247.1719, 238.75, 229.0312, 221.6094, 
    222.3203, 249.8281, 257.2031, 264.6719, 267.5469,
  205, 241, 248.2734, 247.1094, 239.6641, 230.1328, 224.6875, 220.4375, 
    249.6328, 260.4453, 268.6172, 267.8594,
  215.2812, 247.7109, 253.125, 251.7422, 243.5, 228.7188, 220.2969, 219.4609, 
    257.2344, 264.5, 270.7734, 273.3594,
  224.6328, 255.7266, 258.5469, 256.6172, 244.3359, 228.6719, 216.6406, 
    216.9688, 259.9062, 271.4531, 276.875, 283.3984,
  246.0625, 265.5234, 264.5859, 260, 246.5234, 228.1641, 211.3828, 215.5391, 
    258.4531, 270.0312, 276.0703, 278.6641,
  231.0234, 261.8984, 264.8672, 260.5547, 246.9844, 227.5234, 209.9922, 
    215.8047, 253.6172, 271.0312, 280.5234, 286.7188,
  236.7031, 264.6172, 266.4062, 262.3125, 248, 228.9141, 211.4453, 215.4922, 
    253.2891, 270.0391, 280.7266, 287.8906,
  239.8594, 267.6953, 268.0703, 262.8359, 250.3828, 227.7031, 208.0625, 
    215.1328, 251.3984, 267.7656, 277.6953, 285.2969,
  196.3125, 236.3672, 243.4062, 239.875, 227.4531, 212.5703, 203.2109, 
    212.5547, 258.4062, 269.2344, 271.9297, 264.5078,
  220.9766, 246.8984, 249.4297, 244.2891, 232.5781, 218.4297, 211.5391, 
    219.9141, 243.1484, 253.7656, 264.4219, 267.4453,
  201.4375, 240.6797, 246.3594, 243.4688, 232.9766, 222.3984, 217.9219, 
    221.9375, 251.2578, 262.0703, 268.6875, 265.3359,
  227.8125, 248.4766, 248.6719, 244.7969, 235.7344, 227.2812, 221.7812, 
    223.3594, 245.7812, 252.3828, 257.9297, 261.6875,
  211.375, 246.4453, 250.4219, 246.7188, 237.4062, 228.4609, 220.7422, 
    220.9922, 244.4766, 255.0703, 264.5156, 269.625,
  209.9531, 247.4531, 252.3984, 249.1406, 238.0547, 226.3125, 218.0469, 
    219.1328, 255.5391, 264.5391, 270.6484, 273.5938,
  235.0156, 258.9922, 259.5, 253.9844, 242.0312, 223.9609, 213.75, 219.4297, 
    254.6641, 267.7266, 273.5547, 278.6094,
  239.4609, 263.5156, 263.4531, 256.75, 243.9453, 224.1953, 211.4141, 
    215.5469, 254.3672, 268.5703, 275.6641, 279.7969,
  237.1328, 265.7031, 266.1406, 260.125, 245.0234, 224.7266, 209.5547, 
    217.2188, 251.1641, 271.25, 280.5156, 285.9375,
  237.1641, 266.1641, 265.5625, 260.5703, 245.9531, 224.9141, 207.0391, 
    215.8906, 249.4531, 267.4219, 277.1797, 287.2891,
  242.3281, 268.6328, 268.8047, 261.7969, 246.2266, 225.0391, 208.3438, 
    217.6328, 251.7969, 268.1641, 277.5625, 285.25,
  200.3672, 242.1484, 244.1641, 237.2734, 222.2656, 209.0547, 204.1875, 214, 
    252.5859, 265.9609, 271.0391, 270.1484,
  227.4375, 249.8281, 247.8672, 240.8516, 225.9922, 214.8984, 212.2031, 
    219.5781, 237.8203, 249.2188, 260.2344, 267.6016,
  211.6719, 246.2266, 246.4297, 241.0781, 229.7891, 220.1484, 219.0156, 
    223.5469, 240.3672, 253.6406, 263.4922, 267.9375,
  211.1719, 244.8359, 246.1953, 240.5391, 230.9844, 223.5938, 221.0703, 
    222.9453, 237.7891, 246.8125, 255.0703, 262.4453,
  207.6797, 246.5703, 248.9688, 243.3203, 233.9062, 224.9219, 220.1484, 
    222.3281, 245.3438, 256.1172, 265.5312, 270.9766,
  203.6953, 247.4844, 251.375, 246.875, 234.5469, 222.3516, 216.5312, 
    220.6562, 248.6406, 261.6328, 269.7578, 275.375,
  230.5312, 259.5547, 258.8281, 250.3203, 235.5078, 221.6016, 212.2812, 
    219.9375, 250.7031, 266.6172, 272.9922, 279.25,
  244.4297, 264.8281, 261.1562, 252.2422, 237, 219.5156, 209.3906, 219.2812, 
    252.6719, 267.7734, 274.3438, 279.1641,
  245.4922, 269.2266, 265.2656, 254.875, 238.6562, 219.9844, 206.9766, 
    219.1719, 249.5156, 268.7344, 278.6328, 286.0078,
  244.3516, 268.7188, 264.9766, 256.4531, 239.4141, 219.5938, 206.4375, 
    219.9062, 246.6953, 264.3984, 276.1562, 284.8984,
  253.4922, 272.4219, 266.9844, 256.1641, 239.0625, 218.9609, 207.3984, 
    216.7422, 246.5156, 266.5469, 275.2031, 283.0703,
  206.3047, 243.2188, 236.1172, 225.9688, 212.6094, 203.7422, 203.9375, 
    215.5547, 233.5078, 252.3125, 265.0156, 268.0391,
  210.7734, 244.4141, 240.0703, 229.8516, 218.3359, 211.8516, 211.1719, 
    218.5625, 233.0078, 245.6016, 257.4375, 264.1016,
  215.4141, 246.3516, 241.8594, 231.8359, 221.4219, 217.3203, 217.9062, 
    222.7734, 229.9688, 245.3594, 260.3359, 266.8906,
  221.1172, 248.2969, 242.4844, 233.3516, 225.5078, 220.8125, 220.5, 
    224.7344, 240.4141, 251.5156, 262.1328, 268.3984,
  227.0938, 251.0391, 245.875, 236.0938, 226.75, 220.6328, 219.0234, 
    223.5938, 239.6172, 252.1406, 261.8047, 267.9453,
  218.9297, 253.3359, 248.5938, 237.875, 224.4766, 216.9141, 215.7188, 
    222.8047, 234.375, 252.6562, 264.7578, 272.8828,
  240.7656, 261.7578, 253.7578, 241.6953, 226.1172, 215.6562, 214.3672, 
    222.8438, 243.4844, 261.3516, 270.4219, 276.3281,
  259.4609, 265.1484, 255.2188, 242.5391, 225.0703, 213.1406, 210.1172, 
    222.1641, 245.4062, 264.4766, 271.5156, 277.4219,
  262.7969, 269.0078, 258.6406, 245.2109, 227.6875, 212.0859, 207.7969, 
    223.1875, 248.7812, 266.8594, 276.5547, 282.7656,
  273.7344, 269.3438, 259.2344, 244.5312, 226.2656, 212.0859, 206.7734, 
    221.9375, 238.7734, 257.6562, 270.8359, 279.4219,
  264.5781, 269.4531, 259.4922, 245.2031, 227.25, 210.5, 205.7031, 222.5781, 
    236.0234, 259.2969, 269.7734, 280.4453 ;

 clear_fraction =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.3466797, 0.3808594, 0.2900391, 0.3681641, 0.3730469, 0.3720703, 0.375, 
    0.375, 0.3457031, 0.2402344, 0.4033203, 0.4033203,
  0.04003906, 0.03613281, 0.04003906, 0.03710938, 0.03613281, 0.03710938, 
    0.03613281, 0.03613281, 0.07421875, 0.08691406, 0.07128906, 0.07128906,
  0.1679688, 0.1474609, 0.1640625, 0.1523438, 0.1464844, 0.1464844, 
    0.1464844, 0.1464844, 0.1757812, 0.171875, 0.1777344, 0.1767578,
  0.2128906, 0.1757812, 0.1923828, 0.1816406, 0.1816406, 0.1826172, 
    0.1796875, 0.1796875, 0.1552734, 0.1367188, 0.1650391, 0.1640625,
  0.7226562, 0.7539062, 0.7402344, 0.7490234, 0.75, 0.75, 0.7509766, 
    0.7509766, 0.7636719, 0.7822266, 0.7548828, 0.7578125,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.1845703, 0.1582031, 0.171875, 0.1650391, 0.1650391, 0.1650391, 0.1650391, 
    0.1650391, 0.09082031, 0.09765625, 0.078125, 0.078125,
  0.06738281, 0.05566406, 0.05664062, 0.05761719, 0.05761719, 0.05761719, 
    0.05761719, 0.05761719, 0.01171875, 0.01074219, 0.009765625, 0.008789062,
  0.7089844, 0.7041016, 0.7080078, 0.7060547, 0.7060547, 0.7060547, 
    0.7070312, 0.7070312, 0.6757812, 0.6748047, 0.6757812, 0.6767578,
  0.01660156, 0.009765625, 0.01269531, 0.01171875, 0.01171875, 0.01171875, 
    0.01171875, 0.01171875, 0.001953125, 0.001953125, 0.0009765625, 
    0.001953125,
  0.8964844, 0.8974609, 0.8984375, 0.8974609, 0.8964844, 0.8964844, 
    0.8955078, 0.8955078, 0.9199219, 0.9160156, 0.9267578, 0.9257812,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9648438, 0.9609375, 0.9628906, 0.9628906, 0.9628906, 0.9628906, 
    0.9619141, 0.9619141, 0.9707031, 0.9726562, 0.9716797, 0.9716797,
  0.109375, 0.1054688, 0.1083984, 0.1044922, 0.1054688, 0.1054688, 0.1064453, 
    0.1064453, 0.1142578, 0.1142578, 0.1113281, 0.1142578,
  0.7050781, 0.7324219, 0.7216797, 0.7275391, 0.7255859, 0.7246094, 
    0.7255859, 0.7255859, 0.7949219, 0.796875, 0.7958984, 0.796875,
  0.02734375, 0.01757812, 0.02246094, 0.02148438, 0.01953125, 0.01855469, 
    0.01953125, 0.02050781, 0.002929688, 0.002929688, 0.002929688, 0.002929688,
  0.6640625, 0.6953125, 0.6845703, 0.6914062, 0.6904297, 0.6914062, 
    0.6923828, 0.6914062, 0.7207031, 0.7216797, 0.7246094, 0.7246094,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.01953125, 0.006835938, 0.01074219, 0.0078125, 0.008789062, 0.008789062, 
    0.008789062, 0.008789062, 0.001953125, 0.001953125, 0.0009765625, 
    0.0009765625,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.002929688, 0.0009765625, 0.0009765625, 0.0009765625, 0.0009765625, 
    0.0009765625, 0.0009765625, 0.0009765625, 0, 0, 0, 0,
  0.1005859, 0.08007812, 0.0859375, 0.08203125, 0.08203125, 0.08203125, 
    0.08203125, 0.08203125, 0.04589844, 0.04589844, 0.04101562, 0.04003906,
  0.8740234, 0.8828125, 0.8837891, 0.8828125, 0.8818359, 0.8818359, 
    0.8818359, 0.8818359, 0.9492188, 0.9501953, 0.9550781, 0.9560547,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.4648438, 0.4472656, 0.4570312, 0.4521484, 0.4511719, 0.4501953, 
    0.4521484, 0.4521484, 0.4492188, 0.4511719, 0.4326172, 0.4375,
  0.3720703, 0.3876953, 0.3847656, 0.3886719, 0.3847656, 0.3828125, 
    0.3857422, 0.3857422, 0.4042969, 0.40625, 0.4111328, 0.4091797,
  0.2626953, 0.2519531, 0.25, 0.2519531, 0.2548828, 0.2568359, 0.2558594, 
    0.2539062, 0.1621094, 0.1542969, 0.15625, 0.1611328,
  0.5488281, 0.5136719, 0.5234375, 0.5195312, 0.5195312, 0.5195312, 
    0.5175781, 0.5175781, 0.3798828, 0.3769531, 0.3681641, 0.3662109,
  0.6542969, 0.6308594, 0.6347656, 0.6337891, 0.6367188, 0.6376953, 
    0.6367188, 0.6357422, 0.5693359, 0.5664062, 0.5644531, 0.5664062,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0390625, 0.02832031, 0.03320312, 0.02929688, 0.03027344, 0.03027344, 
    0.03027344, 0.03027344, 0.009765625, 0.01074219, 0.005859375, 0.005859375,
  0.6904297, 0.6728516, 0.6767578, 0.6757812, 0.6767578, 0.6777344, 
    0.6787109, 0.6777344, 0.5878906, 0.5859375, 0.5869141, 0.5878906,
  0.8935547, 0.8828125, 0.8876953, 0.8847656, 0.8828125, 0.8828125, 
    0.8837891, 0.8837891, 0.8867188, 0.8886719, 0.8798828, 0.8818359,
  0.890625, 0.9013672, 0.9013672, 0.9003906, 0.9003906, 0.9013672, 0.9013672, 
    0.9013672, 0.9326172, 0.9316406, 0.9355469, 0.9355469,
  0.9462891, 0.9638672, 0.9609375, 0.9619141, 0.9619141, 0.9619141, 
    0.9619141, 0.9619141, 0.984375, 0.9853516, 0.9882812, 0.9882812,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.01269531, 0.002929688, 0.004882812, 0.00390625, 0.00390625, 0.00390625, 
    0.00390625, 0.00390625, 0.001953125, 0.002929688, 0.0009765625, 
    0.0009765625,
  0.08886719, 0.04980469, 0.06347656, 0.05566406, 0.0546875, 0.05566406, 
    0.05566406, 0.05566406, 0.01757812, 0.01953125, 0.0078125, 0.01269531,
  0.8125, 0.8164062, 0.8154297, 0.8164062, 0.8164062, 0.8164062, 0.8173828, 
    0.8173828, 0.8095703, 0.8085938, 0.8164062, 0.8164062,
  0.9912109, 0.9970703, 0.9951172, 0.9960938, 0.9960938, 0.9960938, 
    0.9960938, 0.9960938, 0.9990234, 0.9980469, 0.9990234, 1,
  0.8193359, 0.8330078, 0.8251953, 0.828125, 0.8300781, 0.8300781, 0.828125, 
    0.8271484, 0.9160156, 0.9189453, 0.9257812, 0.9228516,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.7207031, 0.75, 0.7392578, 0.7451172, 0.7431641, 0.7421875, 0.7451172, 
    0.7451172, 0.7548828, 0.7548828, 0.7587891, 0.7587891,
  0.1425781, 0.1279297, 0.1240234, 0.1279297, 0.1289062, 0.1298828, 
    0.1289062, 0.1279297, 0.06445312, 0.05957031, 0.05957031, 0.05761719,
  0.9873047, 0.9931641, 0.9931641, 0.9931641, 0.9931641, 0.9931641, 
    0.9931641, 0.9931641, 0.9990234, 0.9990234, 0.9990234, 1,
  0.8242188, 0.8203125, 0.8222656, 0.8212891, 0.8232422, 0.8232422, 
    0.8212891, 0.8212891, 0.8203125, 0.8164062, 0.8212891, 0.8232422,
  0.9541016, 0.9707031, 0.9638672, 0.9677734, 0.9677734, 0.9677734, 
    0.9667969, 0.9667969, 0.9931641, 0.9931641, 0.9960938, 0.9951172,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.5205078, 0.5058594, 0.5097656, 0.5058594, 0.5097656, 0.5107422, 
    0.5078125, 0.5078125, 0.5576172, 0.5595703, 0.5664062, 0.5664062,
  0.4628906, 0.4736328, 0.4697266, 0.4736328, 0.4707031, 0.46875, 0.4726562, 
    0.4726562, 0.3671875, 0.3603516, 0.3525391, 0.3496094,
  0.6308594, 0.6787109, 0.65625, 0.6689453, 0.6708984, 0.671875, 0.6708984, 
    0.6699219, 0.7636719, 0.7587891, 0.7724609, 0.7734375,
  0.9580078, 0.9628906, 0.9609375, 0.9619141, 0.9628906, 0.9628906, 
    0.9599609, 0.9599609, 0.9970703, 0.9970703, 0.9980469, 0.9980469,
  0.9921875, 0.9941406, 0.9931641, 0.9941406, 0.9951172, 0.9951172, 
    0.9941406, 0.9941406, 0.9990234, 0.9990234, 0.9990234, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.53125, 0.4990234, 0.5136719, 0.5068359, 0.5058594, 0.5058594, 0.5058594, 
    0.5058594, 0.4091797, 0.40625, 0.4003906, 0.3974609,
  0.7041016, 0.6845703, 0.6923828, 0.6894531, 0.6884766, 0.6894531, 
    0.6894531, 0.6894531, 0.6171875, 0.6142578, 0.6123047, 0.6103516,
  0.7226562, 0.7109375, 0.7089844, 0.7109375, 0.7119141, 0.7128906, 
    0.7099609, 0.7099609, 0.6962891, 0.6962891, 0.6982422, 0.6972656,
  0.8701172, 0.890625, 0.8847656, 0.8876953, 0.8867188, 0.8867188, 0.8876953, 
    0.8876953, 0.9257812, 0.9257812, 0.9335938, 0.9326172,
  0.6464844, 0.6474609, 0.6503906, 0.6474609, 0.6464844, 0.6464844, 
    0.6484375, 0.6494141, 0.6650391, 0.6708984, 0.671875, 0.6708984,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.7841797, 0.8066406, 0.8007812, 0.8027344, 0.8037109, 0.8037109, 
    0.8046875, 0.8046875, 0.8476562, 0.8515625, 0.8486328, 0.8515625,
  0.5195312, 0.5488281, 0.5351562, 0.5439453, 0.5429688, 0.5419922, 
    0.5439453, 0.5439453, 0.5595703, 0.5585938, 0.5634766, 0.5625,
  0.859375, 0.8701172, 0.8710938, 0.8671875, 0.8642578, 0.8652344, 0.8671875, 
    0.8671875, 0.9042969, 0.8984375, 0.9140625, 0.9111328,
  0.8730469, 0.8574219, 0.8662109, 0.8603516, 0.859375, 0.859375, 0.8583984, 
    0.8583984, 0.8486328, 0.8544922, 0.8466797, 0.8466797,
  0.9628906, 0.9775391, 0.9726562, 0.9755859, 0.9755859, 0.9755859, 
    0.9765625, 0.9765625, 0.9941406, 0.9951172, 0.9951172, 0.9951172 ;

 cold_target_counts =
  -132995.6, 5.269516e+10, 2.768288e+10, 8.836168e+10, 6.328356e+10, 
    6.934617e+10, 1.649212e+10, 1.836628e+10, -397442, -303380.6, -245941.8, 
    -364101.1,
  -132053.3, 5.284101e+10, 2.774807e+10, 8.854322e+10, 6.340744e+10, 
    6.944133e+10, 1.652521e+10, 1.841952e+10, -396073, -302565.9, -245219.9, 
    -362039.5,
  -131150.1, 5.297147e+10, 2.77931e+10, 8.875431e+10, 6.346818e+10, 
    6.955547e+10, 1.653766e+10, 1.845458e+10, -394799.7, -301371.8, 
    -244338.3, -360133.6,
  -130278.5, 5.312399e+10, 2.783629e+10, 8.882029e+10, 6.354661e+10, 
    6.96589e+10, 1.658267e+10, 1.847216e+10, -394220.8, -301353.6, -243808.5, 
    -359854.7,
  -129248.7, 5.324396e+10, 2.789652e+10, 8.897849e+10, 6.363492e+10, 
    6.973483e+10, 1.658471e+10, 1.8487e+10, -392572.3, -300504.6, -243000.2, 
    -358629.6,
  -128518.4, 5.333777e+10, 2.79165e+10, 8.902033e+10, 6.364501e+10, 
    6.976632e+10, 1.660904e+10, 1.850486e+10, -392175.8, -299748.8, 
    -242314.5, -356876.8,
  -127461.3, 5.350608e+10, 2.798214e+10, 8.926092e+10, 6.381097e+10, 
    6.988829e+10, 1.662746e+10, 1.853291e+10, -391130.3, -299127.2, 
    -241623.6, -356123.2,
  -126775.8, 5.352602e+10, 2.795872e+10, 8.920134e+10, 6.372833e+10, 
    6.985757e+10, 1.661707e+10, 1.851114e+10, -390471.5, -298602.8, 
    -241195.1, -354707.7,
  -125945.9, 5.3645e+10, 2.800392e+10, 8.930304e+10, 6.382658e+10, 
    6.995684e+10, 1.663716e+10, 1.855729e+10, -389345.6, -298256.1, 
    -240659.6, -353671,
  -125297.5, 5.379455e+10, 2.807143e+10, 8.950515e+10, 6.397238e+10, 
    7.008861e+10, 1.667431e+10, 1.860044e+10, -387941.5, -297589.7, 
    -240104.1, -352090.6,
  -124615.7, 5.387599e+10, 2.809942e+10, 8.955494e+10, 6.401267e+10, 
    7.016339e+10, 1.669252e+10, 1.859119e+10, -387596.2, -297512.9, 
    -239418.4, -350918 ;

 combinedQualityFlag =
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1538, 1538, 1538, 1538, 1538, 1538, 1538, 1536, 1536, 1536, 1536,
  1600, 1792, 1536, 1536, 1792, 1536, 1536, 1536, 1920, 1536, 1600, 1808,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536,
  1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1536, 1552,
  1538, 1538, 1538, 1538, 1538, 1538, 1538, 1538, 1538, 1538, 1538, 1554,
  1538, 1538, 1538, 1538, 1538, 1538, 1538, 1538, 1536, 1536, 1536, 1536 ;

 elevation =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1.8125, 0.8125, 0.9375, 0.875, 0.875, 0.875, 0.9375, 0.9375, 0.5, 0.5, 
    0.4375, 0.5,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.125, 0.8125, 0.75, 0.8125, 0.75, 0.75, 0.75, 0.75, 0.3125, 0.3125, 
    0.3125, 0.3125,
  0.0625, 0.0625, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  38.25, 34.5, 33.25, 34.625, 35.3125, 35.5625, 35.125, 34.875, 12.875, 
    12.5625, 11.5625, 11.0625,
  0.3125, 0.1875, 0.125, 0.1875, 0.125, 0.1875, 0.1875, 0.1875, 0.0625, 
    0.0625, 0.0625, 0 ;

 flagAscDesc =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagColdCal =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagDayNight =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 flagICTCal =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagICT_ND_Consistency =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagLunarIntrusion =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagManeuver =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagNDCal =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagNonOcean =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0 ;

 flagOutlierTimestamp =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagPLOrientation =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 flagRFI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagSDRTX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 flagSolarIntrusion =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 instrTemp =
  6.829041, 6.58252, 6.500336, 6.253815, 6.007263, 5.760742, 5.589142, 
    5.424866, 5.26767, 5.103302, 4.946014,
  3.29541, 3.137512, 2.884521, 2.638, 2.562103, 2.309265, 2.144928, 1.892334, 
    1.734039, 1.651886, 1.493408,
  14.40063, 13.82343, 13.14282, 12.51755, 11.92789, 11.25, 10.68918, 10.1221, 
    9.548004, 8.987854, 8.529785,
  14.49994, 13.9032, 13.20303, 12.63898, 12.00949, 11.37384, 10.73096, 
    10.10098, 9.569397, 9.009583, 8.529785,
  14.51981, 13.88324, 13.24316, 12.53781, 11.92789, 11.22931, 10.58472, 
    10.0163, 9.35495, 8.90097, 8.331757,
  14.20187, 13.58371, 13.08246, 12.49731, 11.88696, 11.22931, 10.66837, 
    10.05869, 9.569397, 8.987854, 8.463928 ;

 internal_cal_target_counts =
  -191745.3, 8.587638e+10, 4.4823e+10, 1.51283e+11, 1.085816e+11, 
    1.184951e+11, 2.82814e+10, 3.137509e+10, -536824.2, -399145.3, -339200.6, 
    -472675.8,
  -190545, 8.609871e+10, 4.487747e+10, 1.514054e+11, 1.087131e+11, 
    1.186667e+11, 2.831852e+10, 3.141161e+10, -534678.4, -398007.4, 
    -337940.6, -470357.5,
  -189152.6, 8.633603e+10, 4.497272e+10, 1.516697e+11, 1.089425e+11, 
    1.187233e+11, 2.834702e+10, 3.144374e+10, -533523.1, -396604.7, 
    -336992.4, -468403.9,
  -187966.4, 8.649676e+10, 4.501972e+10, 1.51911e+11, 1.089984e+11, 
    1.188352e+11, 2.838233e+10, 3.147486e+10, -532362.6, -396474.6, 
    -336022.6, -467546.8,
  -186343.3, 8.661886e+10, 4.502817e+10, 1.519118e+11, 1.089913e+11, 
    1.188649e+11, 2.83805e+10, 3.147077e+10, -529911.5, -394750, -334746.1, 
    -465312.5,
  -185056.5, 8.67976e+10, 4.504434e+10, 1.519606e+11, 1.090461e+11, 
    1.189076e+11, 2.840632e+10, 3.150594e+10, -529332.3, -394384.1, 
    -333939.5, -463555.2,
  -183765.5, 8.689608e+10, 4.51495e+10, 1.521529e+11, 1.091407e+11, 
    1.189629e+11, 2.841755e+10, 3.149977e+10, -528209.2, -393435.4, 
    -333093.7, -461925.1,
  -182694.2, 8.697693e+10, 4.510416e+10, 1.520192e+11, 1.090137e+11, 
    1.189232e+11, 2.839934e+10, 3.149279e+10, -526835.7, -392392.7, 
    -332084.4, -460481.7,
  -181536.3, 8.721113e+10, 4.518764e+10, 1.522154e+11, 1.091791e+11, 
    1.191516e+11, 2.842112e+10, 3.155155e+10, -525463.5, -391704, -331335.5, 
    -458878.4,
  -180336.3, 8.734455e+10, 4.526338e+10, 1.524378e+11, 1.092358e+11, 
    1.191711e+11, 2.844068e+10, 3.156543e+10, -523259.8, -391047.7, 
    -330421.9, -456829.2,
  -179285.7, 8.739934e+10, 4.520735e+10, 1.522462e+11, 1.091827e+11, 
    1.19087e+11, 2.844005e+10, 3.153098e+10, -522945.3, -390942.5, -329576, 
    -455427.2 ;

 land_fraction =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.01855469, 0.01660156, 0.01757812, 0.01757812, 0.01757812, 0.01757812, 
    0.01757812, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2724609, 0.2626953, 0.2539062, 0.2626953, 0.265625, 0.2666016, 0.2646484, 
    0.2636719, 0.1679688, 0.1611328, 0.1611328, 0.1591797,
  0.005859375, 0.002929688, 0.002929688, 0.002929688, 0.001953125, 
    0.002929688, 0.002929688, 0.002929688, 0.0009765625, 0.0009765625, 
    0.0009765625, 0 ;

 latitude =
  -50.79004, -45.94629, -41.31738, -36.52051, -31.69629, -26.85449, 
    -21.89648, -16.98535, -12.05371, -7.077148, -2.072266,
  -52.18164, -47.30859, -42.48047, -37.57715, -32.64648, -27.69434, 
    -22.69336, -17.69629, -12.68359, -7.651367, -2.602539,
  -52.77539, -47.86523, -42.96777, -38.01953, -33.04785, -28.05762, 
    -23.03516, -18.00977, -12.97266, -7.920898, -2.858398,
  -53.13477, -48.19824, -43.26172, -38.28711, -33.29297, -28.2832, -23.24805, 
    -18.20801, -13.1582, -8.097656, -3.02832,
  -53.39551, -48.43652, -43.47461, -38.48242, -33.47363, -28.4502, -23.40625, 
    -18.35742, -13.2998, -8.235352, -3.162109,
  -53.6084, -48.63184, -43.65039, -38.64355, -33.62305, -28.59082, -23.54102, 
    -18.48535, -13.42285, -8.355469, -3.28125,
  -53.7998, -48.80762, -43.81055, -38.79102, -33.76172, -28.72168, -23.66699, 
    -18.60742, -13.54199, -8.472656, -3.397461,
  -53.98828, -48.98047, -43.96973, -38.93945, -33.90234, -28.85742, 
    -23.79883, -18.73633, -13.66992, -8.599609, -3.526367,
  -54.18848, -49.16406, -44.14258, -39.10449, -34.06152, -29.0127, -23.95117, 
    -18.88867, -13.82227, -8.755859, -3.68457,
  -54.4043, -49.37109, -44.34473, -39.30176, -34.25781, -29.21094, -24.15137, 
    -19.09277, -14.0332, -8.976562, -3.913086,
  -54.5498, -49.57324, -44.56641, -39.5459, -34.52344, -29.50195, -24.46387, 
    -19.42871, -14.39746, -9.379883, -4.342773 ;

 longitude =
  -0.1621094, -2.678711, -5.670898, -7.861328, -9.854492, -11.74219, 
    -13.03516, -14.55273, -15.9834, -17.16992, -18.1748,
  -5.928711, -8.407227, -10.84473, -12.79004, -14.53223, -16.13086, 
    -17.43066, -18.75, -19.98535, -21.10352, -22.12207,
  -8.986328, -11.30176, -13.47754, -15.26367, -16.8623, -18.33008, -19.58203, 
    -20.81445, -21.97754, -23.06055, -24.07129,
  -11.12793, -13.28613, -15.2832, -16.95117, -18.44824, -19.82715, -21.0332, 
    -22.20801, -23.32812, -24.38672, -25.38965,
  -12.875, -14.88184, -16.73438, -18.30078, -19.71875, -21.02637, -22.18945, 
    -23.31738, -24.40332, -25.44434, -26.43945,
  -14.47266, -16.32227, -18.04492, -19.51465, -20.86035, -22.10449, 
    -23.22461, -24.31348, -25.36719, -26.3916, -27.37988,
  -16.08496, -17.76074, -19.35449, -20.72363, -21.99219, -23.17676, -24.25, 
    -25.30273, -26.32617, -27.33301, -28.3125,
  -17.89648, -19.34961, -20.80664, -22.05859, -23.24023, -24.36035, 
    -25.37695, -26.39258, -27.38477, -28.37109, -29.33789,
  -20.19043, -21.32324, -22.61816, -23.7207, -24.79297, -25.83398, -26.77441, 
    -27.74121, -28.69531, -29.66309, -30.60938,
  -23.60938, -24.18652, -25.25781, -26.13379, -27.04785, -27.97852, 
    -28.79883, -29.68652, -30.58984, -31.54004, -32.44727,
  -30.53613, -29.66797, -30.36523, -30.76758, -31.38184, -32.125, -32.67285, 
    -33.37891, -34.19043, -35.15625, -35.96289 ;

 lunar_azimuth_angle =
  71.14062, 70.75781, 70.59375, 69.75781, 68.71875, 67.55469, 66.14844, 
    64.82812, 63.50781, 62.20312, 60.97656,
  75.78906, 74.98438, 74.02344, 72.60938, 71.00781, 69.29688, 67.46875, 
    65.69531, 63.95312, 62.28125, 60.71875,
  78.29688, 77.16406, 75.78906, 74.05469, 72.15625, 70.16406, 68.10938, 
    66.10156, 64.15625, 62.29688, 60.5625,
  80.07031, 78.66406, 77.01562, 75.04688, 72.92969, 70.75, 68.53125, 
    66.36719, 64.28125, 62.29688, 60.44531,
  81.51562, 79.875, 78, 75.84375, 73.55469, 71.21875, 68.86719, 66.57812, 
    64.375, 62.28906, 60.34375,
  82.85156, 80.97656, 78.89062, 76.55469, 74.11719, 71.64062, 69.16406, 
    66.75781, 64.45312, 62.28125, 60.25,
  84.20312, 82.07812, 79.78125, 77.26562, 74.67188, 72.05469, 69.45312, 
    66.9375, 64.53125, 62.26562, 60.14844,
  85.72656, 83.29688, 80.77344, 78.05469, 75.28125, 72.50781, 69.76562, 
    67.125, 64.60938, 62.24219, 60.03125,
  87.66406, 84.82031, 82.02344, 79.03906, 76.04688, 73.07031, 70.14844, 
    67.35156, 64.69531, 62.20312, 59.875,
  90.57031, 87.04688, 83.83594, 80.46875, 77.14062, 73.88281, 70.69531, 
    67.66406, 64.80469, 62.125, 59.63281,
  96.52344, 91.32812, 87.36719, 83.20312, 79.22656, 75.40625, 71.67969, 
    68.20312, 64.94531, 61.90625, 59.10156 ;

 lunar_zenith_angle =
  112.8281, 112.625, 112.9141, 112.6641, 112.25, 111.7188, 110.5938, 
    109.5859, 108.4141, 106.9141, 105.1406,
  116.6328, 116.7578, 116.9062, 116.6953, 116.2656, 115.6328, 114.6172, 
    113.5, 112.1719, 110.6094, 108.8203,
  118.5703, 118.7656, 118.8906, 118.6797, 118.2344, 117.5625, 116.5703, 
    115.4062, 114.0391, 112.4375, 110.6328,
  119.8906, 120.125, 120.2266, 120.0156, 119.5625, 118.875, 117.875, 
    116.6875, 115.2891, 113.6719, 111.8516,
  120.9531, 121.2031, 121.2969, 121.0859, 120.625, 119.9141, 118.9141, 
    117.7109, 116.2891, 114.6562, 112.8281,
  121.9141, 122.1641, 122.25, 122.0312, 121.5703, 120.8516, 119.8438, 
    118.6172, 117.1797, 115.5391, 113.6953,
  122.875, 123.1172, 123.2031, 122.9766, 122.5078, 121.7734, 120.7578, 
    119.5234, 118.0625, 116.4141, 114.5547,
  123.9453, 124.1719, 124.25, 124.0156, 123.5312, 122.7969, 121.7578, 
    120.5156, 119.0391, 117.3672, 115.5,
  125.2891, 125.4609, 125.5469, 125.2969, 124.8047, 124.0625, 123, 121.7344, 
    120.25, 118.5625, 116.6641,
  127.2656, 127.3203, 127.4297, 127.1562, 126.6484, 125.8984, 124.7891, 
    123.5, 121.9844, 120.2891, 118.3516,
  131.2266, 130.8438, 131.0469, 130.6953, 130.1641, 129.4219, 128.2031, 
    126.8203, 125.2656, 123.6016, 121.5625 ;

 noise_diode_counts =
  -189247.3, 8.040816e+10, 4.066503e+10, 1.35206e+11, 9.715824e+10, 
    1.060862e+11, 2.509706e+10, 2.770851e+10, -538287.3, -387948.3, 
    -354664.3, -446341.2,
  -188321.3, 8.07584e+10, 4.077033e+10, 1.355951e+11, 9.742779e+10, 
    1.063825e+11, 2.517703e+10, 2.781688e+10, -537089.4, -387101.4, 
    -353648.3, -444513.3,
  -187141.3, 8.095774e+10, 4.084595e+10, 1.359355e+11, 9.755243e+10, 
    1.06537e+11, 2.518675e+10, 2.78376e+10, -536294.9, -386092, -352909.3, 
    -442719.2,
  -185985.8, 8.112506e+10, 4.087995e+10, 1.360508e+11, 9.759933e+10, 
    1.066135e+11, 2.523457e+10, 2.789349e+10, -535123.6, -385670.1, 
    -352248.3, -441870.1,
  -184525.7, 8.140951e+10, 4.09984e+10, 1.363596e+11, 9.781997e+10, 
    1.067936e+11, 2.526175e+10, 2.790641e+10, -532790.6, -384562.9, 
    -351163.9, -440137.8,
  -183509.8, 8.168634e+10, 4.105949e+10, 1.36521e+11, 9.796959e+10, 
    1.069674e+11, 2.531632e+10, 2.795033e+10, -532805.1, -384418.8, 
    -350619.1, -439038.7,
  -182274.5, 8.18459e+10, 4.116104e+10, 1.368383e+11, 9.820516e+10, 
    1.071e+11, 2.532848e+10, 2.799948e+10, -531840.6, -383370.7, -349788.2, 
    -437482.4,
  -181282.1, 8.20445e+10, 4.122014e+10, 1.369971e+11, 9.828139e+10, 
    1.072021e+11, 2.537763e+10, 2.800975e+10, -530938.5, -382833.1, 
    -349089.7, -436080.2,
  -180277.5, 8.227926e+10, 4.129862e+10, 1.372525e+11, 9.842634e+10, 
    1.074478e+11, 2.543184e+10, 2.809744e+10, -529951.1, -382788.9, 
    -348821.2, -435337.1,
  -179535.4, 8.244003e+10, 4.138194e+10, 1.374326e+11, 9.851692e+10, 
    1.07543e+11, 2.546194e+10, 2.813215e+10, -528291.2, -382050.6, -348049.7, 
    -433336.7,
  -178653.5, 8.260229e+10, 4.138739e+10, 1.37534e+11, 9.860482e+10, 
    1.076668e+11, 2.547179e+10, 2.817047e+10, -527984.5, -381950.6, 
    -347258.2, -431595.2 ;

 scAltitude = 508.363, 506.488, 504.5078, 502.467, 500.4279, 498.4368, 
    496.5409, 494.792, 493.2231, 491.8722, 490.7614 ;

 scLatitude = -53.56514, -48.60619, -43.62116, -38.6164, -33.5956, -28.56149, 
    -23.51643, -18.46238, -13.40096, -8.333833, -3.263057 ;

 scLongitude = -14.41477, -16.40089, -18.09196, -19.57568, -20.91004, 
    -22.13493, -23.27908, -24.36394, -25.40629, -26.41985, -27.41626 ;

 scPosECEF =
  3969.17, -1020.2, -5517.141,
  4374.733, -1287.627, -5141.673,
  4743.136, -1549.559, -4725.77,
  5071.498, -1803.454, -4272.725,
  5357.349, -2046.848, -3786.072,
  5598.567, -2277.32, -3269.607,
  5793.392, -2492.521, -2727.39,
  5940.466, -2690.208, -2163.685,
  6038.827, -2868.259, -1582.903,
  6087.919, -3024.698, -989.6185,
  6087.592, -3157.7, -388.5534 ;

 scQuatECEF =
  0.1917415, 0.3313575, 0.07313422, -0.9209174,
  0.1913154, 0.3724246, 0.06322408, -0.9059255,
  0.1896147, 0.4121431, 0.05075537, -0.8897237,
  0.1872339, 0.451063, 0.03799119, -0.8718041,
  0.1844538, 0.4890161, 0.02484351, -0.8521871,
  0.1812128, 0.5259356, 0.01148894, -0.8309162,
  0.1774956, 0.5617562, -0.002125079, -0.8080351,
  0.1732616, 0.5964037, -0.01592017, -0.7836004,
  0.1685978, 0.6297906, -0.02992402, -0.7576563,
  0.1634, 0.6619213, -0.04400208, -0.7302222,
  0.15776, 0.6926353, -0.05824269, -0.7014099 ;

 scRollAngle = 10.05804, 10.01935, 10.00567, 10.01904, 10.01898, 10.00936, 
    10.00607, 10.02268, 10.03029, 10.01315, 10.01578 ;

 scVelECEF =
  5.289881, -3.367281, 4.428906,
  4.843697, -3.313857, 4.952698,
  4.360273, -3.229079, 5.437954,
  3.843642, -3.113136, 5.880902,
  3.298207, -2.966623, 6.277656,
  2.728578, -2.790246, 6.62535,
  2.139257, -2.585068, 6.921138,
  1.535517, -2.352646, 7.162426,
  0.9222055, -2.094488, 7.347376,
  0.3045877, -1.812646, 7.474526,
  -0.3123069, -1.509181, 7.542591 ;

 sensor_azimuth_angle =
  246.7334, 248.9902, 251.6514, 253.665, 255.4326, 257.0186, 258.2383, 
    259.4668, 260.5586, 261.5059, 262.3662,
  251.3789, 253.2891, 255.2412, 256.7676, 258.0547, 259.1572, 260.0254, 
    260.8311, 261.5195, 262.1055, 262.6113,
  254.0059, 255.626, 257.2285, 258.4824, 259.5127, 260.375, 261.04, 261.6318, 
    262.1172, 262.5146, 262.833,
  256.0957, 257.4668, 258.833, 259.8867, 260.7383, 261.4316, 261.9375, 
    262.374, 262.7109, 262.9668, 263.1387,
  258.625, 259.6699, 260.8613, 261.7314, 262.4336, 262.9863, 263.3008, 
    263.5771, 263.7617, 263.8701, 263.8623,
  38.59863, 296.2646, 310.4297, 299.5859, 303.7627, 317.2686, 296.1826, 
    295.3018, 300.2354, 307.748, 296.3057,
  77.10938, 77.64062, 78.51465, 79.0918, 79.61328, 80.07617, 80.3623, 
    80.66211, 80.92578, 81.11426, 81.24512,
  79.56641, 80.00391, 80.65039, 81.08105, 81.43066, 81.70605, 81.86426, 
    81.99609, 82.07324, 82.08594, 82.05078,
  81.7832, 81.88965, 82.29883, 82.51855, 82.68164, 82.78516, 82.78516, 
    82.76367, 82.69043, 82.56152, 82.38477,
  84.75391, 84.27051, 84.34863, 84.25195, 84.15332, 84.02441, 83.7998, 
    83.57422, 83.30957, 83.00098, 82.64062,
  90.52344, 88.57715, 88.06445, 87.33203, 86.7373, 86.1875, 85.51953, 
    84.9082, 84.30078, 83.67676, 82.98242 ;

 sensor_view_angle =
  59.87402, 60.89355, 60.56152, 60.77246, 60.82422, 60.64648, 61.13379, 
    60.98242, 60.73438, 60.7207, 60.87012,
  47.78223, 48.83008, 48.51172, 48.72266, 48.75391, 48.5752, 49.03125, 
    48.8877, 48.67676, 48.64941, 48.80176,
  35.69824, 36.76562, 36.45117, 36.65723, 36.69238, 36.49609, 36.92188, 
    36.78906, 36.59082, 36.55273, 36.71582,
  23.61426, 24.69824, 24.39551, 24.59277, 24.62109, 24.41309, 24.80273, 
    24.7002, 24.50781, 24.44824, 24.61426,
  11.53223, 12.63184, 12.36719, 12.55176, 12.53125, 12.33398, 12.67871, 
    12.62988, 12.46191, 12.3623, 12.50781,
  -0.6884766, 0.7294922, 0.5683594, 0.6962891, 0.6376953, 0.5058594, 
    0.7089844, 0.6884766, 0.5664062, 0.4521484, 0.5205078,
  -12.55371, -11.4248, -11.61426, -11.42285, -11.50586, -11.69531, -11.42188, 
    -11.44727, -11.53613, -11.66016, -11.57324,
  -24.55273, -23.37402, -23.56934, -23.36328, -23.43359, -23.63965, 
    -23.37891, -23.44238, -23.50293, -23.62305, -23.54395,
  -36.56836, -35.29785, -35.54199, -35.33301, -35.39062, -35.60449, 
    -35.34766, -35.42383, -35.47852, -35.62695, -35.52441,
  -48.56738, -47.20312, -47.50684, -47.30762, -47.36133, -47.57617, 
    -47.32422, -47.36621, -47.42969, -47.63965, -47.50195,
  -60.52148, -59.09668, -59.44043, -59.26074, -59.32129, -59.53125, 
    -59.29297, -59.25195, -59.32715, -59.62109, -59.45703 ;

 sensor_zenith_angle =
  69.02441, 70.55957, 69.99805, 70.28223, 70.31836, 70, 70.71875, 70.44141, 
    70.02148, 69.9707, 70.17578,
  53.08398, 54.33496, 53.92676, 54.16016, 54.17676, 53.93848, 54.47168, 
    54.27832, 54.00488, 53.95703, 54.12793,
  39.04492, 40.24023, 39.87109, 40.09082, 40.11719, 39.88281, 40.35156, 
    40.19043, 39.95605, 39.90332, 40.0791,
  25.62207, 26.80566, 26.46582, 26.67383, 26.69629, 26.46094, 26.88086, 
    26.76172, 26.54492, 26.47363, 26.65039,
  12.46387, 13.65137, 13.36133, 13.55762, 13.53125, 13.31445, 13.68359, 
    13.62793, 13.44238, 13.33203, 13.48828,
  0.7431641, 0.7871094, 0.6132812, 0.7509766, 0.6884766, 0.5449219, 
    0.7646484, 0.7421875, 0.609375, 0.4873047, 0.5615234,
  13.57031, 12.34473, 12.5459, 12.33594, 12.42188, 12.62305, 12.32422, 
    12.34961, 12.44141, 12.57422, 12.47754,
  26.65234, 25.35156, 25.55859, 25.32617, 25.39551, 25.61328, 25.32031, 
    25.38379, 25.44434, 25.57031, 25.47949,
  40.02832, 38.58105, 38.84375, 38.59668, 38.64844, 38.87793, 38.57617, 
    38.65137, 38.70215, 38.86035, 38.73828,
  54.0332, 52.36621, 52.71094, 52.45117, 52.49512, 52.73242, 52.41113, 
    52.44434, 52.50391, 52.74121, 52.56445,
  70.01367, 67.82617, 68.2959, 67.99121, 68.04102, 68.3125, 67.9248, 
    67.83105, 67.91016, 68.31445, 68.05176 ;

 solar_azimuth_angle =
  171.1016, 173.5078, 177.1328, 180.1328, 183.6016, 188.0781, 192.9062, 
    201.4688, 216.0547, 241.3516, 276.7344,
  178.8672, 181.8438, 185.3203, 188.7578, 192.7891, 197.875, 204.2891, 
    213.8125, 227.9688, 248.1641, 272.1797,
  182.875, 185.9141, 189.3203, 192.875, 197.0703, 202.3516, 209.125, 
    218.7031, 232.2188, 250.2969, 270.9297,
  185.6406, 188.6484, 192, 195.5938, 199.8672, 205.2344, 212.1406, 221.6562, 
    234.6719, 251.4766, 270.2969,
  187.875, 190.8203, 194.125, 197.7266, 202.0391, 207.4609, 214.4141, 
    223.8203, 236.4219, 252.3125, 269.875,
  189.8984, 192.7578, 196.0078, 199.6094, 203.9531, 209.3906, 216.3516, 
    225.6406, 237.8594, 252.9922, 269.5469,
  191.9219, 194.6719, 197.8672, 201.4531, 205.7969, 211.25, 218.1875, 
    227.3438, 239.1797, 253.6094, 269.2656,
  194.1719, 196.7656, 199.9062, 203.4453, 207.7891, 213.2344, 220.125, 
    229.1094, 240.5312, 254.2422, 268.9922,
  197, 199.3359, 202.3984, 205.8828, 210.1875, 215.6094, 222.3984, 231.1484, 
    242.0703, 254.9531, 268.7031,
  201.1562, 203, 205.9609, 209.3125, 213.5469, 218.8984, 225.4688, 233.8359, 
    244.0625, 255.8828, 268.3594,
  209.3828, 209.8125, 212.5859, 215.5781, 219.5938, 224.7188, 230.7344, 
    238.2891, 247.2969, 257.4219, 267.9062 ;

 solar_beta_angle = 18.76284, 18.80257, 18.78373, 18.70697, 18.57521, 
    18.39212, 18.16399, 17.8981, 17.60276, 17.28737, 16.96194 ;

 solar_zenith_angle =
  131.8906, 136.8828, 141.6562, 146.4844, 151.2578, 155.9375, 160.6562, 
    165.0312, 168.875, 171.5938, 171.8984,
  130.8203, 135.6797, 140.4062, 145.125, 149.75, 154.2422, 158.6016, 
    162.5312, 165.7734, 167.8125, 168.0078,
  130.1953, 134.9922, 139.6797, 144.3203, 148.8594, 153.2344, 157.4062, 
    161.1172, 164.1016, 165.9062, 166.0703,
  129.7422, 134.4922, 139.1406, 143.7344, 148.2109, 152.4922, 156.5391, 
    160.1094, 162.9297, 164.6094, 164.75,
  129.3594, 134.0781, 138.6953, 143.2422, 147.6562, 151.875, 155.8281, 
    159.2812, 161.9922, 163.5703, 163.7031,
  129, 133.6953, 138.2812, 142.7891, 147.1484, 151.3047, 155.1641, 158.5312, 
    161.1328, 162.6406, 162.7656,
  128.6328, 133.2969, 137.8516, 142.3203, 146.625, 150.7109, 154.4922, 
    157.7656, 160.2734, 161.7109, 161.8359,
  128.2109, 132.8516, 137.3672, 141.7812, 146.0312, 150.0469, 153.7422, 
    156.9062, 159.3281, 160.6953, 160.8125,
  127.6562, 132.2734, 136.7344, 141.0938, 145.2734, 149.1875, 152.7891, 
    155.8359, 158.1328, 159.4219, 159.5391,
  126.7969, 131.4062, 135.7734, 140.0547, 144.1172, 147.8984, 151.3594, 
    154.25, 156.3984, 157.5703, 157.6953,
  124.9531, 129.6406, 133.7969, 137.9297, 141.7734, 145.2656, 148.5234, 
    151.1719, 153.0703, 154, 154.1797 ;
}
